module shifter(out, shamt, left, sign, in);
	output [63:0] out;
	input [5:0] shamt;
	input left, sign;
	input [63:0] in;
	
	wire invLeft, top;
	wire [6:0] sel, invSel;
	wire [63:-3] stage1;
	wire [63:-15] stage2;
	wire [63:-63] stage3;
	
	//selection logic
	and SE(top, sign, in[63]);
	xor x5(sel[5], shamt[5], left);
	xor x4(sel[4], shamt[4], left);
	xor x3(sel[3], shamt[3], left);
	xor x2(sel[2], shamt[2], left);
	xor x1(sel[1], shamt[1], left);
	xor x0(sel[0], shamt[0], left);
	not n5(invSel[5], sel[5]);
	not n4(invSel[4], sel[4]);
	not n3(invSel[3], sel[3]);
	not n2(invSel[2], sel[2]);
	not n1(invSel[1], sel[1]);
	not n0(invSel[0], sel[0]);
	not nL(invLeft, left);
	
	//first stage, 63--3
		NAND_MUX_4x1 mux0_neg3(.out(stage1[-3]), .select(sel[1:0]), .invSelect(invSel[1:0]), .in({in[0], 3'h0}));
	NAND_MUX_4x1 mux0_neg2(.out(stage1[-2]), .select(sel[1:0]), .invSelect(invSel[1:0]), .in({in[1:0], 2'h0}));
	NAND_MUX_4x1 mux0_neg1(.out(stage1[-1]), .select(sel[1:0]), .invSelect(invSel[1:0]), .in({in[2:0], 1'b0}));
	//NAND_MUX_4x1 mux0_neg0(.out(stage1[-0], .select(sel[1:0]), .invSelect(invSel[1:0]), .in({in3:0]));
		NAND_MUX_4x1 mux0_7(.out(stage1[7]), .select(sel[1:0]), .invSelect(invSel[1:0]), .in(in[10:7]));
	NAND_MUX_4x1 mux0_6(.out(stage1[6]), .select(sel[1:0]), .invSelect(invSel[1:0]), .in(in[9:6]));
	NAND_MUX_4x1 mux0_5(.out(stage1[5]), .select(sel[1:0]), .invSelect(invSel[1:0]), .in(in[8:5]));
	NAND_MUX_4x1 mux0_4(.out(stage1[4]), .select(sel[1:0]), .invSelect(invSel[1:0]), .in(in[7:4]));
	NAND_MUX_4x1 mux0_3(.out(stage1[3]), .select(sel[1:0]), .invSelect(invSel[1:0]), .in(in[6:3]));
	NAND_MUX_4x1 mux0_2(.out(stage1[2]), .select(sel[1:0]), .invSelect(invSel[1:0]), .in(in[5:2]));
	NAND_MUX_4x1 mux0_1(.out(stage1[1]), .select(sel[1:0]), .invSelect(invSel[1:0]), .in(in[4:1]));
	NAND_MUX_4x1 mux0_0(.out(stage1[0]), .select(sel[1:0]), .invSelect(invSel[1:0]), .in(in[3:0]));
		NAND_MUX_4x1 mux0_15(.out(stage1[15]), .select(sel[1:0]), .invSelect(invSel[1:0]), .in(in[18:15]));
	NAND_MUX_4x1 mux0_14(.out(stage1[14]), .select(sel[1:0]), .invSelect(invSel[1:0]), .in(in[17:14]));
	NAND_MUX_4x1 mux0_13(.out(stage1[13]), .select(sel[1:0]), .invSelect(invSel[1:0]), .in(in[16:13]));
	NAND_MUX_4x1 mux0_12(.out(stage1[12]), .select(sel[1:0]), .invSelect(invSel[1:0]), .in(in[15:12]));
	NAND_MUX_4x1 mux0_11(.out(stage1[11]), .select(sel[1:0]), .invSelect(invSel[1:0]), .in(in[14:11]));
	NAND_MUX_4x1 mux0_10(.out(stage1[10]), .select(sel[1:0]), .invSelect(invSel[1:0]), .in(in[13:10]));
	NAND_MUX_4x1 mux0_9(.out(stage1[9]), .select(sel[1:0]), .invSelect(invSel[1:0]), .in(in[12:9]));
	NAND_MUX_4x1 mux0_8(.out(stage1[8]), .select(sel[1:0]), .invSelect(invSel[1:0]), .in(in[11:8]));
		NAND_MUX_4x1 mux0_23(.out(stage1[23]), .select(sel[1:0]), .invSelect(invSel[1:0]), .in(in[26:23]));
	NAND_MUX_4x1 mux0_22(.out(stage1[22]), .select(sel[1:0]), .invSelect(invSel[1:0]), .in(in[25:22]));
	NAND_MUX_4x1 mux0_21(.out(stage1[21]), .select(sel[1:0]), .invSelect(invSel[1:0]), .in(in[24:21]));
	NAND_MUX_4x1 mux0_20(.out(stage1[20]), .select(sel[1:0]), .invSelect(invSel[1:0]), .in(in[23:20]));
	NAND_MUX_4x1 mux0_19(.out(stage1[19]), .select(sel[1:0]), .invSelect(invSel[1:0]), .in(in[22:19]));
	NAND_MUX_4x1 mux0_18(.out(stage1[18]), .select(sel[1:0]), .invSelect(invSel[1:0]), .in(in[21:18]));
	NAND_MUX_4x1 mux0_17(.out(stage1[17]), .select(sel[1:0]), .invSelect(invSel[1:0]), .in(in[20:17]));
	NAND_MUX_4x1 mux0_16(.out(stage1[16]), .select(sel[1:0]), .invSelect(invSel[1:0]), .in(in[19:16]));
		NAND_MUX_4x1 mux0_31(.out(stage1[31]), .select(sel[1:0]), .invSelect(invSel[1:0]), .in(in[34:31]));
	NAND_MUX_4x1 mux0_30(.out(stage1[30]), .select(sel[1:0]), .invSelect(invSel[1:0]), .in(in[33:30]));
	NAND_MUX_4x1 mux0_29(.out(stage1[29]), .select(sel[1:0]), .invSelect(invSel[1:0]), .in(in[32:29]));
	NAND_MUX_4x1 mux0_28(.out(stage1[28]), .select(sel[1:0]), .invSelect(invSel[1:0]), .in(in[31:28]));
	NAND_MUX_4x1 mux0_27(.out(stage1[27]), .select(sel[1:0]), .invSelect(invSel[1:0]), .in(in[30:27]));
	NAND_MUX_4x1 mux0_26(.out(stage1[26]), .select(sel[1:0]), .invSelect(invSel[1:0]), .in(in[29:26]));
	NAND_MUX_4x1 mux0_25(.out(stage1[25]), .select(sel[1:0]), .invSelect(invSel[1:0]), .in(in[28:25]));
	NAND_MUX_4x1 mux0_24(.out(stage1[24]), .select(sel[1:0]), .invSelect(invSel[1:0]), .in(in[27:24]));
		NAND_MUX_4x1 mux0_39(.out(stage1[39]), .select(sel[1:0]), .invSelect(invSel[1:0]), .in(in[42:39]));
	NAND_MUX_4x1 mux0_38(.out(stage1[38]), .select(sel[1:0]), .invSelect(invSel[1:0]), .in(in[41:38]));
	NAND_MUX_4x1 mux0_37(.out(stage1[37]), .select(sel[1:0]), .invSelect(invSel[1:0]), .in(in[40:37]));
	NAND_MUX_4x1 mux0_36(.out(stage1[36]), .select(sel[1:0]), .invSelect(invSel[1:0]), .in(in[39:36]));
	NAND_MUX_4x1 mux0_35(.out(stage1[35]), .select(sel[1:0]), .invSelect(invSel[1:0]), .in(in[38:35]));
	NAND_MUX_4x1 mux0_34(.out(stage1[34]), .select(sel[1:0]), .invSelect(invSel[1:0]), .in(in[37:34]));
	NAND_MUX_4x1 mux0_33(.out(stage1[33]), .select(sel[1:0]), .invSelect(invSel[1:0]), .in(in[36:33]));
	NAND_MUX_4x1 mux0_32(.out(stage1[32]), .select(sel[1:0]), .invSelect(invSel[1:0]), .in(in[35:32]));
		NAND_MUX_4x1 mux0_47(.out(stage1[47]), .select(sel[1:0]), .invSelect(invSel[1:0]), .in(in[50:47]));
	NAND_MUX_4x1 mux0_46(.out(stage1[46]), .select(sel[1:0]), .invSelect(invSel[1:0]), .in(in[49:46]));
	NAND_MUX_4x1 mux0_45(.out(stage1[45]), .select(sel[1:0]), .invSelect(invSel[1:0]), .in(in[48:45]));
	NAND_MUX_4x1 mux0_44(.out(stage1[44]), .select(sel[1:0]), .invSelect(invSel[1:0]), .in(in[47:44]));
	NAND_MUX_4x1 mux0_43(.out(stage1[43]), .select(sel[1:0]), .invSelect(invSel[1:0]), .in(in[46:43]));
	NAND_MUX_4x1 mux0_42(.out(stage1[42]), .select(sel[1:0]), .invSelect(invSel[1:0]), .in(in[45:42]));
	NAND_MUX_4x1 mux0_41(.out(stage1[41]), .select(sel[1:0]), .invSelect(invSel[1:0]), .in(in[44:41]));
	NAND_MUX_4x1 mux0_40(.out(stage1[40]), .select(sel[1:0]), .invSelect(invSel[1:0]), .in(in[43:40]));
		NAND_MUX_4x1 mux0_55(.out(stage1[55]), .select(sel[1:0]), .invSelect(invSel[1:0]), .in(in[58:55]));
	NAND_MUX_4x1 mux0_54(.out(stage1[54]), .select(sel[1:0]), .invSelect(invSel[1:0]), .in(in[57:54]));
	NAND_MUX_4x1 mux0_53(.out(stage1[53]), .select(sel[1:0]), .invSelect(invSel[1:0]), .in(in[56:53]));
	NAND_MUX_4x1 mux0_52(.out(stage1[52]), .select(sel[1:0]), .invSelect(invSel[1:0]), .in(in[55:52]));
	NAND_MUX_4x1 mux0_51(.out(stage1[51]), .select(sel[1:0]), .invSelect(invSel[1:0]), .in(in[54:51]));
	NAND_MUX_4x1 mux0_50(.out(stage1[50]), .select(sel[1:0]), .invSelect(invSel[1:0]), .in(in[53:50]));
	NAND_MUX_4x1 mux0_49(.out(stage1[49]), .select(sel[1:0]), .invSelect(invSel[1:0]), .in(in[52:49]));
	NAND_MUX_4x1 mux0_48(.out(stage1[48]), .select(sel[1:0]), .invSelect(invSel[1:0]), .in(in[51:48]));
		NAND_MUX_4x1 mux0_63(.out(stage1[63]), .select(sel[1:0]), .invSelect(invSel[1:0]), .in({{3{top}}, in[63]}));
	NAND_MUX_4x1 mux0_62(.out(stage1[62]), .select(sel[1:0]), .invSelect(invSel[1:0]), .in({{2{top}}, in[63:62]}));
	NAND_MUX_4x1 mux0_61(.out(stage1[61]), .select(sel[1:0]), .invSelect(invSel[1:0]), .in({top, in[63:61]}));
	NAND_MUX_4x1 mux0_60(.out(stage1[60]), .select(sel[1:0]), .invSelect(invSel[1:0]), .in(in[63:60]));
	NAND_MUX_4x1 mux0_59(.out(stage1[59]), .select(sel[1:0]), .invSelect(invSel[1:0]), .in(in[62:59]));
	NAND_MUX_4x1 mux0_58(.out(stage1[58]), .select(sel[1:0]), .invSelect(invSel[1:0]), .in(in[61:58]));
	NAND_MUX_4x1 mux0_57(.out(stage1[57]), .select(sel[1:0]), .invSelect(invSel[1:0]), .in(in[60:57]));
	NAND_MUX_4x1 mux0_56(.out(stage1[56]), .select(sel[1:0]), .invSelect(invSel[1:0]), .in(in[59:56]));
	
	//second stage, 63--15
		NAND_MUX_4x1 mux1_neg15(.out(stage2[-15]), .select(sel[3:2]), .invSelect(invSel[3:2]), .in({stage1[-3], 3'h0}));
	NAND_MUX_4x1 mux1_neg14(.out(stage2[-14]), .select(sel[3:2]), .invSelect(invSel[3:2]), .in({stage1[-2], 3'h0}));
	NAND_MUX_4x1 mux1_neg13(.out(stage2[-13]), .select(sel[3:2]), .invSelect(invSel[3:2]), .in({stage1[-1], 3'h0}));
	NAND_MUX_4x1 mux1_neg12(.out(stage2[-12]), .select(sel[3:2]), .invSelect(invSel[3:2]), .in({stage1[0], 3'h0}));
	NAND_MUX_4x1 mux1_neg11(.out(stage2[-11]), .select(sel[3:2]), .invSelect(invSel[3:2]), .in({stage1[1], stage1[-3], 2'h0}));
	NAND_MUX_4x1 mux1_neg10(.out(stage2[-10]), .select(sel[3:2]), .invSelect(invSel[3:2]), .in({stage1[2], stage1[-2], 2'h0}));
	NAND_MUX_4x1 mux1_neg9(.out(stage2[-9]), .select(sel[3:2]), .invSelect(invSel[3:2]), .in({stage1[3], stage1[-1], 2'h0}));
	NAND_MUX_4x1 mux1_neg8(.out(stage2[-8]), .select(sel[3:2]), .invSelect(invSel[3:2]), .in({stage1[4], stage1[0], 2'h0}));
		NAND_MUX_4x1 mux1_neg7(.out(stage2[-7]), .select(sel[3:2]), .invSelect(invSel[3:2]), .in({stage1[5], stage1[1], stage1[-3], 1'b0}));
	NAND_MUX_4x1 mux1_neg6(.out(stage2[-6]), .select(sel[3:2]), .invSelect(invSel[3:2]), .in({stage1[6], stage1[2], stage1[-2], 1'b0}));
	NAND_MUX_4x1 mux1_neg5(.out(stage2[-5]), .select(sel[3:2]), .invSelect(invSel[3:2]), .in({stage1[7], stage1[3], stage1[-1], 1'b0}));
	NAND_MUX_4x1 mux1_neg4(.out(stage2[-4]), .select(sel[3:2]), .invSelect(invSel[3:2]), .in({stage1[8], stage1[4], stage1[0], 1'b0}));
	NAND_MUX_4x1 mux1_neg3(.out(stage2[-3]), .select(sel[3:2]), .invSelect(invSel[3:2]), .in({stage1[9], stage1[5], stage1[1], stage1[-3]}));
	NAND_MUX_4x1 mux1_neg2(.out(stage2[-2]), .select(sel[3:2]), .invSelect(invSel[3:2]), .in({stage1[10], stage1[6], stage1[2], stage1[-2]}));
	NAND_MUX_4x1 mux1_neg1(.out(stage2[-1]), .select(sel[3:2]), .invSelect(invSel[3:2]), .in({stage1[11], stage1[7], stage1[3], stage1[-1]}));
	//NAND_MUX_4x1 mux1_neg0(.out(stage2[-0]), .select(sel[3:2]), .invSelect(invSel[3:2]), .in({stage1[12], stage1[8], stage1[4], stage1[0]}));
		NAND_MUX_4x1 mux1_7(.out(stage2[7]), .select(sel[3:2]), .invSelect(invSel[3:2]), .in({stage1[19], stage1[15], stage1[11], stage1[7]}));
	NAND_MUX_4x1 mux1_6(.out(stage2[6]), .select(sel[3:2]), .invSelect(invSel[3:2]), .in({stage1[18], stage1[14], stage1[10], stage1[6]}));
	NAND_MUX_4x1 mux1_5(.out(stage2[5]), .select(sel[3:2]), .invSelect(invSel[3:2]), .in({stage1[17], stage1[13], stage1[9], stage1[5]}));
	NAND_MUX_4x1 mux1_4(.out(stage2[4]), .select(sel[3:2]), .invSelect(invSel[3:2]), .in({stage1[16], stage1[12], stage1[8], stage1[4]}));
	NAND_MUX_4x1 mux1_3(.out(stage2[3]), .select(sel[3:2]), .invSelect(invSel[3:2]), .in({stage1[15], stage1[11], stage1[7], stage1[3]}));
	NAND_MUX_4x1 mux1_2(.out(stage2[2]), .select(sel[3:2]), .invSelect(invSel[3:2]), .in({stage1[14], stage1[10], stage1[6], stage1[2]}));
	NAND_MUX_4x1 mux1_1(.out(stage2[1]), .select(sel[3:2]), .invSelect(invSel[3:2]), .in({stage1[13], stage1[9], stage1[5], stage1[1]}));
	NAND_MUX_4x1 mux1_0(.out(stage2[0]), .select(sel[3:2]), .invSelect(invSel[3:2]), .in({stage1[12], stage1[8], stage1[4], stage1[0]}));
		NAND_MUX_4x1 mux1_15(.out(stage2[15]), .select(sel[3:2]), .invSelect(invSel[3:2]), .in({stage1[27], stage1[23], stage1[19], stage1[15]}));
	NAND_MUX_4x1 mux1_14(.out(stage2[14]), .select(sel[3:2]), .invSelect(invSel[3:2]), .in({stage1[26], stage1[22], stage1[18], stage1[14]}));
	NAND_MUX_4x1 mux1_13(.out(stage2[13]), .select(sel[3:2]), .invSelect(invSel[3:2]), .in({stage1[25], stage1[21], stage1[17], stage1[13]}));
	NAND_MUX_4x1 mux1_12(.out(stage2[12]), .select(sel[3:2]), .invSelect(invSel[3:2]), .in({stage1[24], stage1[20], stage1[16], stage1[12]}));
	NAND_MUX_4x1 mux1_11(.out(stage2[11]), .select(sel[3:2]), .invSelect(invSel[3:2]), .in({stage1[23], stage1[19], stage1[15], stage1[11]}));
	NAND_MUX_4x1 mux1_10(.out(stage2[10]), .select(sel[3:2]), .invSelect(invSel[3:2]), .in({stage1[22], stage1[18], stage1[14], stage1[10]}));
	NAND_MUX_4x1 mux1_9(.out(stage2[9]), .select(sel[3:2]), .invSelect(invSel[3:2]), .in({stage1[21], stage1[17], stage1[13], stage1[9]}));
	NAND_MUX_4x1 mux1_8(.out(stage2[8]), .select(sel[3:2]), .invSelect(invSel[3:2]), .in({stage1[20], stage1[16], stage1[12], stage1[8]}));
		NAND_MUX_4x1 mux1_23(.out(stage2[23]), .select(sel[3:2]), .invSelect(invSel[3:2]), .in({stage1[35], stage1[31], stage1[27], stage1[23]}));
	NAND_MUX_4x1 mux1_22(.out(stage2[22]), .select(sel[3:2]), .invSelect(invSel[3:2]), .in({stage1[34], stage1[30], stage1[26], stage1[22]}));
	NAND_MUX_4x1 mux1_21(.out(stage2[21]), .select(sel[3:2]), .invSelect(invSel[3:2]), .in({stage1[33], stage1[29], stage1[25], stage1[21]}));
	NAND_MUX_4x1 mux1_20(.out(stage2[20]), .select(sel[3:2]), .invSelect(invSel[3:2]), .in({stage1[32], stage1[28], stage1[24], stage1[20]}));
	NAND_MUX_4x1 mux1_19(.out(stage2[19]), .select(sel[3:2]), .invSelect(invSel[3:2]), .in({stage1[31], stage1[27], stage1[23], stage1[19]}));
	NAND_MUX_4x1 mux1_18(.out(stage2[18]), .select(sel[3:2]), .invSelect(invSel[3:2]), .in({stage1[30], stage1[26], stage1[22], stage1[18]}));
	NAND_MUX_4x1 mux1_17(.out(stage2[17]), .select(sel[3:2]), .invSelect(invSel[3:2]), .in({stage1[29], stage1[25], stage1[21], stage1[17]}));
	NAND_MUX_4x1 mux1_16(.out(stage2[16]), .select(sel[3:2]), .invSelect(invSel[3:2]), .in({stage1[28], stage1[24], stage1[20], stage1[16]}));
		NAND_MUX_4x1 mux1_31(.out(stage2[31]), .select(sel[3:2]), .invSelect(invSel[3:2]), .in({stage1[43], stage1[39], stage1[35], stage1[31]}));
	NAND_MUX_4x1 mux1_30(.out(stage2[30]), .select(sel[3:2]), .invSelect(invSel[3:2]), .in({stage1[42], stage1[38], stage1[34], stage1[30]}));
	NAND_MUX_4x1 mux1_29(.out(stage2[29]), .select(sel[3:2]), .invSelect(invSel[3:2]), .in({stage1[41], stage1[37], stage1[33], stage1[29]}));
	NAND_MUX_4x1 mux1_28(.out(stage2[28]), .select(sel[3:2]), .invSelect(invSel[3:2]), .in({stage1[40], stage1[36], stage1[32], stage1[28]}));
	NAND_MUX_4x1 mux1_27(.out(stage2[27]), .select(sel[3:2]), .invSelect(invSel[3:2]), .in({stage1[39], stage1[35], stage1[31], stage1[27]}));
	NAND_MUX_4x1 mux1_26(.out(stage2[26]), .select(sel[3:2]), .invSelect(invSel[3:2]), .in({stage1[38], stage1[34], stage1[30], stage1[26]}));
	NAND_MUX_4x1 mux1_25(.out(stage2[25]), .select(sel[3:2]), .invSelect(invSel[3:2]), .in({stage1[37], stage1[33], stage1[29], stage1[25]}));
	NAND_MUX_4x1 mux1_24(.out(stage2[24]), .select(sel[3:2]), .invSelect(invSel[3:2]), .in({stage1[36], stage1[32], stage1[28], stage1[24]}));
		NAND_MUX_4x1 mux1_39(.out(stage2[39]), .select(sel[3:2]), .invSelect(invSel[3:2]), .in({stage1[51], stage1[47], stage1[43], stage1[39]}));
	NAND_MUX_4x1 mux1_38(.out(stage2[38]), .select(sel[3:2]), .invSelect(invSel[3:2]), .in({stage1[50], stage1[46], stage1[42], stage1[38]}));
	NAND_MUX_4x1 mux1_37(.out(stage2[37]), .select(sel[3:2]), .invSelect(invSel[3:2]), .in({stage1[49], stage1[45], stage1[41], stage1[37]}));
	NAND_MUX_4x1 mux1_36(.out(stage2[36]), .select(sel[3:2]), .invSelect(invSel[3:2]), .in({stage1[48], stage1[44], stage1[40], stage1[36]}));
	NAND_MUX_4x1 mux1_35(.out(stage2[35]), .select(sel[3:2]), .invSelect(invSel[3:2]), .in({stage1[47], stage1[43], stage1[39], stage1[35]}));
	NAND_MUX_4x1 mux1_34(.out(stage2[34]), .select(sel[3:2]), .invSelect(invSel[3:2]), .in({stage1[46], stage1[42], stage1[38], stage1[34]}));
	NAND_MUX_4x1 mux1_33(.out(stage2[33]), .select(sel[3:2]), .invSelect(invSel[3:2]), .in({stage1[45], stage1[41], stage1[37], stage1[33]}));
	NAND_MUX_4x1 mux1_32(.out(stage2[32]), .select(sel[3:2]), .invSelect(invSel[3:2]), .in({stage1[44], stage1[40], stage1[36], stage1[32]}));
		NAND_MUX_4x1 mux1_47(.out(stage2[47]), .select(sel[3:2]), .invSelect(invSel[3:2]), .in({stage1[59], stage1[55], stage1[51], stage1[47]}));
	NAND_MUX_4x1 mux1_46(.out(stage2[46]), .select(sel[3:2]), .invSelect(invSel[3:2]), .in({stage1[58], stage1[54], stage1[50], stage1[46]}));
	NAND_MUX_4x1 mux1_45(.out(stage2[45]), .select(sel[3:2]), .invSelect(invSel[3:2]), .in({stage1[57], stage1[53], stage1[49], stage1[45]}));
	NAND_MUX_4x1 mux1_44(.out(stage2[44]), .select(sel[3:2]), .invSelect(invSel[3:2]), .in({stage1[56], stage1[52], stage1[48], stage1[44]}));
	NAND_MUX_4x1 mux1_43(.out(stage2[43]), .select(sel[3:2]), .invSelect(invSel[3:2]), .in({stage1[55], stage1[51], stage1[47], stage1[43]}));
	NAND_MUX_4x1 mux1_42(.out(stage2[42]), .select(sel[3:2]), .invSelect(invSel[3:2]), .in({stage1[54], stage1[50], stage1[46], stage1[42]}));
	NAND_MUX_4x1 mux1_41(.out(stage2[41]), .select(sel[3:2]), .invSelect(invSel[3:2]), .in({stage1[53], stage1[49], stage1[45], stage1[41]}));
	NAND_MUX_4x1 mux1_40(.out(stage2[40]), .select(sel[3:2]), .invSelect(invSel[3:2]), .in({stage1[52], stage1[48], stage1[44], stage1[40]}));
		NAND_MUX_4x1 mux1_55(.out(stage2[55]), .select(sel[3:2]), .invSelect(invSel[3:2]), .in({top, stage1[63], stage1[59], stage1[55]}));
	NAND_MUX_4x1 mux1_54(.out(stage2[54]), .select(sel[3:2]), .invSelect(invSel[3:2]), .in({top, stage1[62], stage1[58], stage1[54]}));
	NAND_MUX_4x1 mux1_53(.out(stage2[53]), .select(sel[3:2]), .invSelect(invSel[3:2]), .in({top, stage1[61], stage1[57], stage1[53]}));
	NAND_MUX_4x1 mux1_52(.out(stage2[52]), .select(sel[3:2]), .invSelect(invSel[3:2]), .in({top, stage1[60], stage1[56], stage1[52]}));
	NAND_MUX_4x1 mux1_51(.out(stage2[51]), .select(sel[3:2]), .invSelect(invSel[3:2]), .in({stage1[63], stage1[59], stage1[55], stage1[51]}));
	NAND_MUX_4x1 mux1_50(.out(stage2[50]), .select(sel[3:2]), .invSelect(invSel[3:2]), .in({stage1[62], stage1[58], stage1[54], stage1[50]}));
	NAND_MUX_4x1 mux1_49(.out(stage2[49]), .select(sel[3:2]), .invSelect(invSel[3:2]), .in({stage1[61], stage1[57], stage1[53], stage1[49]}));
	NAND_MUX_4x1 mux1_48(.out(stage2[48]), .select(sel[3:2]), .invSelect(invSel[3:2]), .in({stage1[60], stage1[56], stage1[52], stage1[48]}));
		NAND_MUX_4x1 mux1_63(.out(stage2[63]), .select(sel[3:2]), .invSelect(invSel[3:2]), .in({{3{top}}, stage1[63]}));
	NAND_MUX_4x1 mux1_62(.out(stage2[62]), .select(sel[3:2]), .invSelect(invSel[3:2]), .in({{3{top}}, stage1[62]}));
	NAND_MUX_4x1 mux1_61(.out(stage2[61]), .select(sel[3:2]), .invSelect(invSel[3:2]), .in({{3{top}}, stage1[61]}));
	NAND_MUX_4x1 mux1_60(.out(stage2[60]), .select(sel[3:2]), .invSelect(invSel[3:2]), .in({{3{top}}, stage1[60]}));
	NAND_MUX_4x1 mux1_59(.out(stage2[59]), .select(sel[3:2]), .invSelect(invSel[3:2]), .in({{2{top}}, stage1[63], stage1[59]}));
	NAND_MUX_4x1 mux1_58(.out(stage2[58]), .select(sel[3:2]), .invSelect(invSel[3:2]), .in({{2{top}}, stage1[62], stage1[58]}));
	NAND_MUX_4x1 mux1_57(.out(stage2[57]), .select(sel[3:2]), .invSelect(invSel[3:2]), .in({{2{top}}, stage1[61], stage1[57]}));
	NAND_MUX_4x1 mux1_56(.out(stage2[56]), .select(sel[3:2]), .invSelect(invSel[3:2]), .in({{2{top}}, stage1[60], stage1[56]}));
	
	//stage 3, shift 63--63
		NAND_MUX_4x1 mux2_neg63(.out(stage3[-63]), .select(sel[5:4]), .invSelect(invSel[5:4]), .in({stage2[-15], 3'h0}));
	NAND_MUX_4x1 mux2_neg62(.out(stage3[-62]), .select(sel[5:4]), .invSelect(invSel[5:4]), .in({stage2[-14], 3'h0}));
	NAND_MUX_4x1 mux2_neg61(.out(stage3[-61]), .select(sel[5:4]), .invSelect(invSel[5:4]), .in({stage2[-13], 3'h0}));
	NAND_MUX_4x1 mux2_neg60(.out(stage3[-60]), .select(sel[5:4]), .invSelect(invSel[5:4]), .in({stage2[-12], 3'h0}));
	NAND_MUX_4x1 mux2_neg59(.out(stage3[-59]), .select(sel[5:4]), .invSelect(invSel[5:4]), .in({stage2[-11], 3'h0}));
	NAND_MUX_4x1 mux2_neg58(.out(stage3[-58]), .select(sel[5:4]), .invSelect(invSel[5:4]), .in({stage2[-10], 3'h0}));
	NAND_MUX_4x1 mux2_neg57(.out(stage3[-57]), .select(sel[5:4]), .invSelect(invSel[5:4]), .in({stage2[-9], 3'h0}));
	NAND_MUX_4x1 mux2_neg56(.out(stage3[-56]), .select(sel[5:4]), .invSelect(invSel[5:4]), .in({stage2[-8], 3'h0}));
		NAND_MUX_4x1 mux2_neg55(.out(stage3[-55]), .select(sel[5:4]), .invSelect(invSel[5:4]), .in({stage2[-7], 3'h0}));
	NAND_MUX_4x1 mux2_neg54(.out(stage3[-54]), .select(sel[5:4]), .invSelect(invSel[5:4]), .in({stage2[-6], 3'h0}));
	NAND_MUX_4x1 mux2_neg53(.out(stage3[-53]), .select(sel[5:4]), .invSelect(invSel[5:4]), .in({stage2[-5], 3'h0}));
	NAND_MUX_4x1 mux2_neg52(.out(stage3[-52]), .select(sel[5:4]), .invSelect(invSel[5:4]), .in({stage2[-4], 3'h0}));
	NAND_MUX_4x1 mux2_neg51(.out(stage3[-51]), .select(sel[5:4]), .invSelect(invSel[5:4]), .in({stage2[-3], 3'h0}));
	NAND_MUX_4x1 mux2_neg50(.out(stage3[-50]), .select(sel[5:4]), .invSelect(invSel[5:4]), .in({stage2[-2], 3'h0}));
	NAND_MUX_4x1 mux2_neg49(.out(stage3[-49]), .select(sel[5:4]), .invSelect(invSel[5:4]), .in({stage2[-1], 3'h0}));
	NAND_MUX_4x1 mux2_neg48(.out(stage3[-48]), .select(sel[5:4]), .invSelect(invSel[5:4]), .in({stage2[0], 3'h0}));
		NAND_MUX_4x1 mux2_neg47(.out(stage3[-47]), .select(sel[5:4]), .invSelect(invSel[5:4]), .in({stage2[1], stage2[-15], 2'h0}));
	NAND_MUX_4x1 mux2_neg46(.out(stage3[-46]), .select(sel[5:4]), .invSelect(invSel[5:4]), .in({stage2[2], stage2[-14], 2'h0}));
	NAND_MUX_4x1 mux2_neg45(.out(stage3[-45]), .select(sel[5:4]), .invSelect(invSel[5:4]), .in({stage2[3], stage2[-13], 2'h0}));
	NAND_MUX_4x1 mux2_neg44(.out(stage3[-44]), .select(sel[5:4]), .invSelect(invSel[5:4]), .in({stage2[4], stage2[-12], 2'h0}));
	NAND_MUX_4x1 mux2_neg43(.out(stage3[-43]), .select(sel[5:4]), .invSelect(invSel[5:4]), .in({stage2[5], stage2[-11], 2'h0}));
	NAND_MUX_4x1 mux2_neg42(.out(stage3[-42]), .select(sel[5:4]), .invSelect(invSel[5:4]), .in({stage2[6], stage2[-10], 2'h0}));
	NAND_MUX_4x1 mux2_neg41(.out(stage3[-41]), .select(sel[5:4]), .invSelect(invSel[5:4]), .in({stage2[7], stage2[-9], 2'h0}));
	NAND_MUX_4x1 mux2_neg40(.out(stage3[-40]), .select(sel[5:4]), .invSelect(invSel[5:4]), .in({stage2[8], stage2[-8], 2'h0}));
		NAND_MUX_4x1 mux2_neg39(.out(stage3[-39]), .select(sel[5:4]), .invSelect(invSel[5:4]), .in({stage2[9], stage2[-7], 2'h0}));
	NAND_MUX_4x1 mux2_neg38(.out(stage3[-38]), .select(sel[5:4]), .invSelect(invSel[5:4]), .in({stage2[10], stage2[-6], 2'h0}));
	NAND_MUX_4x1 mux2_neg37(.out(stage3[-37]), .select(sel[5:4]), .invSelect(invSel[5:4]), .in({stage2[11], stage2[-5], 2'h0}));
	NAND_MUX_4x1 mux2_neg36(.out(stage3[-36]), .select(sel[5:4]), .invSelect(invSel[5:4]), .in({stage2[12], stage2[-4], 2'h0}));
	NAND_MUX_4x1 mux2_neg35(.out(stage3[-35]), .select(sel[5:4]), .invSelect(invSel[5:4]), .in({stage2[13], stage2[-3], 2'h0}));
	NAND_MUX_4x1 mux2_neg34(.out(stage3[-34]), .select(sel[5:4]), .invSelect(invSel[5:4]), .in({stage2[14], stage2[-2], 2'h0}));
	NAND_MUX_4x1 mux2_neg33(.out(stage3[-33]), .select(sel[5:4]), .invSelect(invSel[5:4]), .in({stage2[15], stage2[-1], 2'h0}));
	NAND_MUX_4x1 mux2_neg32(.out(stage3[-32]), .select(sel[5:4]), .invSelect(invSel[5:4]), .in({stage2[16], stage2[0], 2'h0}));
		NAND_MUX_4x1 mux2_neg31(.out(stage3[-31]), .select(sel[5:4]), .invSelect(invSel[5:4]), .in({stage2[17], stage2[1], stage2[-15], 1'h0}));
	NAND_MUX_4x1 mux2_neg30(.out(stage3[-30]), .select(sel[5:4]), .invSelect(invSel[5:4]), .in({stage2[18], stage2[2], stage2[-14], 1'h0}));
	NAND_MUX_4x1 mux2_neg29(.out(stage3[-29]), .select(sel[5:4]), .invSelect(invSel[5:4]), .in({stage2[19], stage2[3], stage2[-13], 1'h0}));
	NAND_MUX_4x1 mux2_neg28(.out(stage3[-28]), .select(sel[5:4]), .invSelect(invSel[5:4]), .in({stage2[20], stage2[4], stage2[-12], 1'h0}));
	NAND_MUX_4x1 mux2_neg27(.out(stage3[-27]), .select(sel[5:4]), .invSelect(invSel[5:4]), .in({stage2[21], stage2[5], stage2[-11], 1'h0}));
	NAND_MUX_4x1 mux2_neg26(.out(stage3[-26]), .select(sel[5:4]), .invSelect(invSel[5:4]), .in({stage2[22], stage2[6], stage2[-10], 1'h0}));
	NAND_MUX_4x1 mux2_neg25(.out(stage3[-25]), .select(sel[5:4]), .invSelect(invSel[5:4]), .in({stage2[23], stage2[7], stage2[-9], 1'h0}));
	NAND_MUX_4x1 mux2_neg24(.out(stage3[-24]), .select(sel[5:4]), .invSelect(invSel[5:4]), .in({stage2[24], stage2[8], stage2[-8], 1'h0}));
		NAND_MUX_4x1 mux2_neg23(.out(stage3[-23]), .select(sel[5:4]), .invSelect(invSel[5:4]), .in({stage2[25], stage2[9], stage2[-7], 1'h0}));
	NAND_MUX_4x1 mux2_neg22(.out(stage3[-22]), .select(sel[5:4]), .invSelect(invSel[5:4]), .in({stage2[26], stage2[10], stage2[-6], 1'h0}));
	NAND_MUX_4x1 mux2_neg21(.out(stage3[-21]), .select(sel[5:4]), .invSelect(invSel[5:4]), .in({stage2[27], stage2[11], stage2[-5], 1'h0}));
	NAND_MUX_4x1 mux2_neg20(.out(stage3[-20]), .select(sel[5:4]), .invSelect(invSel[5:4]), .in({stage2[28], stage2[12], stage2[-4], 1'h0}));
	NAND_MUX_4x1 mux2_neg19(.out(stage3[-19]), .select(sel[5:4]), .invSelect(invSel[5:4]), .in({stage2[29], stage2[13], stage2[-3], 1'h0}));
	NAND_MUX_4x1 mux2_neg18(.out(stage3[-18]), .select(sel[5:4]), .invSelect(invSel[5:4]), .in({stage2[30], stage2[14], stage2[-2], 1'h0}));
	NAND_MUX_4x1 mux2_neg17(.out(stage3[-17]), .select(sel[5:4]), .invSelect(invSel[5:4]), .in({stage2[31], stage2[15], stage2[-1], 1'h0}));
	NAND_MUX_4x1 mux2_neg16(.out(stage3[-16]), .select(sel[5:4]), .invSelect(invSel[5:4]), .in({stage2[32], stage2[16], stage2[0], 1'h0}));
		NAND_MUX_4x1 mux2_neg15(.out(stage3[-15]), .select(sel[5:4]), .invSelect(invSel[5:4]), .in({stage2[33], stage2[17], stage2[1], stage2[-15]}));
	NAND_MUX_4x1 mux2_neg14(.out(stage3[-14]), .select(sel[5:4]), .invSelect(invSel[5:4]), .in({stage2[34], stage2[18], stage2[2], stage2[-14]}));
	NAND_MUX_4x1 mux2_neg13(.out(stage3[-13]), .select(sel[5:4]), .invSelect(invSel[5:4]), .in({stage2[35], stage2[19], stage2[3], stage2[-13]}));
	NAND_MUX_4x1 mux2_neg12(.out(stage3[-12]), .select(sel[5:4]), .invSelect(invSel[5:4]), .in({stage2[36], stage2[20], stage2[4], stage2[-12]}));
	NAND_MUX_4x1 mux2_neg11(.out(stage3[-11]), .select(sel[5:4]), .invSelect(invSel[5:4]), .in({stage2[37], stage2[21], stage2[5], stage2[-11]}));
	NAND_MUX_4x1 mux2_neg10(.out(stage3[-10]), .select(sel[5:4]), .invSelect(invSel[5:4]), .in({stage2[38], stage2[22], stage2[6], stage2[-10]}));
	NAND_MUX_4x1 mux2_neg9(.out(stage3[-9]), .select(sel[5:4]), .invSelect(invSel[5:4]), .in({stage2[39], stage2[23], stage2[7], stage2[-9]}));
	NAND_MUX_4x1 mux2_neg8(.out(stage3[-8]), .select(sel[5:4]), .invSelect(invSel[5:4]), .in({stage2[40], stage2[24], stage2[8], stage2[-8]}));
		NAND_MUX_4x1 mux2_neg7(.out(stage3[-7]), .select(sel[5:4]), .invSelect(invSel[5:4]), .in({stage2[41], stage2[25], stage2[9], stage2[-7]}));
	NAND_MUX_4x1 mux2_neg6(.out(stage3[-6]), .select(sel[5:4]), .invSelect(invSel[5:4]), .in({stage2[42], stage2[26], stage2[10], stage2[-6]}));
	NAND_MUX_4x1 mux2_neg5(.out(stage3[-5]), .select(sel[5:4]), .invSelect(invSel[5:4]), .in({stage2[43], stage2[27], stage2[11], stage2[-5]}));
	NAND_MUX_4x1 mux2_neg4(.out(stage3[-4]), .select(sel[5:4]), .invSelect(invSel[5:4]), .in({stage2[44], stage2[28], stage2[12], stage2[-4]}));
	NAND_MUX_4x1 mux2_neg3(.out(stage3[-3]), .select(sel[5:4]), .invSelect(invSel[5:4]), .in({stage2[45], stage2[29], stage2[13], stage2[-3]}));
	NAND_MUX_4x1 mux2_neg2(.out(stage3[-2]), .select(sel[5:4]), .invSelect(invSel[5:4]), .in({stage2[46], stage2[30], stage2[14], stage2[-2]}));
	NAND_MUX_4x1 mux2_neg1(.out(stage3[-1]), .select(sel[5:4]), .invSelect(invSel[5:4]), .in({stage2[47], stage2[31], stage2[15], stage2[-1]}));
	//NAND_MUX_4x1 mux2_neg0(.out(stage3[-0]), .select(sel[5:4]), .invSelect(invSel[5:4]), .in({stage2[48], stage2[32], stage2[16], stage2[0]}));
		NAND_MUX_4x1 mux2_7(.out(stage3[7]), .select(sel[5:4]), .invSelect(invSel[5:4]), .in({stage2[55], stage2[39], stage2[23], stage2[7]}));
	NAND_MUX_4x1 mux2_6(.out(stage3[6]), .select(sel[5:4]), .invSelect(invSel[5:4]), .in({stage2[54], stage2[38], stage2[22], stage2[6]}));
	NAND_MUX_4x1 mux2_5(.out(stage3[5]), .select(sel[5:4]), .invSelect(invSel[5:4]), .in({stage2[53], stage2[37], stage2[21], stage2[5]}));
	NAND_MUX_4x1 mux2_4(.out(stage3[4]), .select(sel[5:4]), .invSelect(invSel[5:4]), .in({stage2[52], stage2[36], stage2[20], stage2[4]}));
	NAND_MUX_4x1 mux2_3(.out(stage3[3]), .select(sel[5:4]), .invSelect(invSel[5:4]), .in({stage2[51], stage2[35], stage2[19], stage2[3]}));
	NAND_MUX_4x1 mux2_2(.out(stage3[2]), .select(sel[5:4]), .invSelect(invSel[5:4]), .in({stage2[50], stage2[34], stage2[18], stage2[2]}));
	NAND_MUX_4x1 mux2_1(.out(stage3[1]), .select(sel[5:4]), .invSelect(invSel[5:4]), .in({stage2[49], stage2[33], stage2[17], stage2[1]}));
	NAND_MUX_4x1 mux2_0(.out(stage3[0]), .select(sel[5:4]), .invSelect(invSel[5:4]), .in({stage2[48], stage2[32], stage2[16], stage2[0]}));
		NAND_MUX_4x1 mux2_15(.out(stage3[15]), .select(sel[5:4]), .invSelect(invSel[5:4]), .in({stage2[63], stage2[47], stage2[31], stage2[15]}));
	NAND_MUX_4x1 mux2_14(.out(stage3[14]), .select(sel[5:4]), .invSelect(invSel[5:4]), .in({stage2[62], stage2[46], stage2[30], stage2[14]}));
	NAND_MUX_4x1 mux2_13(.out(stage3[13]), .select(sel[5:4]), .invSelect(invSel[5:4]), .in({stage2[61], stage2[45], stage2[29], stage2[13]}));
	NAND_MUX_4x1 mux2_12(.out(stage3[12]), .select(sel[5:4]), .invSelect(invSel[5:4]), .in({stage2[60], stage2[44], stage2[28], stage2[12]}));
	NAND_MUX_4x1 mux2_11(.out(stage3[11]), .select(sel[5:4]), .invSelect(invSel[5:4]), .in({stage2[59], stage2[43], stage2[27], stage2[11]}));
	NAND_MUX_4x1 mux2_10(.out(stage3[10]), .select(sel[5:4]), .invSelect(invSel[5:4]), .in({stage2[58], stage2[42], stage2[26], stage2[10]}));
	NAND_MUX_4x1 mux2_9(.out(stage3[9]), .select(sel[5:4]), .invSelect(invSel[5:4]), .in({stage2[57], stage2[41], stage2[25], stage2[9]}));
	NAND_MUX_4x1 mux2_8(.out(stage3[8]), .select(sel[5:4]), .invSelect(invSel[5:4]), .in({stage2[56], stage2[40], stage2[24], stage2[8]}));
		NAND_MUX_4x1 mux2_23(.out(stage3[23]), .select(sel[5:4]), .invSelect(invSel[5:4]), .in({1'b0, stage2[55], stage2[39], stage2[23]}));
	NAND_MUX_4x1 mux2_22(.out(stage3[22]), .select(sel[5:4]), .invSelect(invSel[5:4]), .in({top, stage2[54], stage2[38], stage2[22]}));
	NAND_MUX_4x1 mux2_21(.out(stage3[21]), .select(sel[5:4]), .invSelect(invSel[5:4]), .in({top, stage2[53], stage2[37], stage2[21]}));
	NAND_MUX_4x1 mux2_20(.out(stage3[20]), .select(sel[5:4]), .invSelect(invSel[5:4]), .in({top, stage2[52], stage2[36], stage2[20]}));
	NAND_MUX_4x1 mux2_19(.out(stage3[19]), .select(sel[5:4]), .invSelect(invSel[5:4]), .in({top, stage2[51], stage2[35], stage2[19]}));
	NAND_MUX_4x1 mux2_18(.out(stage3[18]), .select(sel[5:4]), .invSelect(invSel[5:4]), .in({top, stage2[50], stage2[34], stage2[18]}));
	NAND_MUX_4x1 mux2_17(.out(stage3[17]), .select(sel[5:4]), .invSelect(invSel[5:4]), .in({top, stage2[49], stage2[33], stage2[17]}));
	NAND_MUX_4x1 mux2_16(.out(stage3[16]), .select(sel[5:4]), .invSelect(invSel[5:4]), .in({top, stage2[48], stage2[32], stage2[16]}));
		NAND_MUX_4x1 mux2_31(.out(stage3[31]), .select(sel[5:4]), .invSelect(invSel[5:4]), .in({top, stage2[63], stage2[47], stage2[31]}));
	NAND_MUX_4x1 mux2_30(.out(stage3[30]), .select(sel[5:4]), .invSelect(invSel[5:4]), .in({top, stage2[62], stage2[46], stage2[30]}));
	NAND_MUX_4x1 mux2_29(.out(stage3[29]), .select(sel[5:4]), .invSelect(invSel[5:4]), .in({top, stage2[61], stage2[45], stage2[29]}));
	NAND_MUX_4x1 mux2_28(.out(stage3[28]), .select(sel[5:4]), .invSelect(invSel[5:4]), .in({top, stage2[60], stage2[44], stage2[28]}));
	NAND_MUX_4x1 mux2_27(.out(stage3[27]), .select(sel[5:4]), .invSelect(invSel[5:4]), .in({top, stage2[59], stage2[43], stage2[27]}));
	NAND_MUX_4x1 mux2_26(.out(stage3[26]), .select(sel[5:4]), .invSelect(invSel[5:4]), .in({top, stage2[58], stage2[42], stage2[26]}));
	NAND_MUX_4x1 mux2_25(.out(stage3[25]), .select(sel[5:4]), .invSelect(invSel[5:4]), .in({top, stage2[57], stage2[41], stage2[25]}));
	NAND_MUX_4x1 mux2_24(.out(stage3[24]), .select(sel[5:4]), .invSelect(invSel[5:4]), .in({top, stage2[56], stage2[40], stage2[24]}));
		NAND_MUX_4x1 mux2_39(.out(stage3[39]), .select(sel[5:4]), .invSelect(invSel[5:4]), .in({{2{top}}, stage2[55], stage2[39]}));
	NAND_MUX_4x1 mux2_38(.out(stage3[38]), .select(sel[5:4]), .invSelect(invSel[5:4]), .in({{2{top}}, stage2[54], stage2[38]}));
	NAND_MUX_4x1 mux2_37(.out(stage3[37]), .select(sel[5:4]), .invSelect(invSel[5:4]), .in({{2{top}}, stage2[53], stage2[37]}));
	NAND_MUX_4x1 mux2_36(.out(stage3[36]), .select(sel[5:4]), .invSelect(invSel[5:4]), .in({{2{top}}, stage2[52], stage2[36]}));
	NAND_MUX_4x1 mux2_35(.out(stage3[35]), .select(sel[5:4]), .invSelect(invSel[5:4]), .in({{2{top}}, stage2[51], stage2[35]}));
	NAND_MUX_4x1 mux2_34(.out(stage3[34]), .select(sel[5:4]), .invSelect(invSel[5:4]), .in({{2{top}}, stage2[50], stage2[34]}));
	NAND_MUX_4x1 mux2_33(.out(stage3[33]), .select(sel[5:4]), .invSelect(invSel[5:4]), .in({{2{top}}, stage2[49], stage2[33]}));
	NAND_MUX_4x1 mux2_32(.out(stage3[32]), .select(sel[5:4]), .invSelect(invSel[5:4]), .in({{2{top}}, stage2[48], stage2[32]}));
		NAND_MUX_4x1 mux2_47(.out(stage3[47]), .select(sel[5:4]), .invSelect(invSel[5:4]), .in({{2{top}}, stage2[63], stage2[47]}));
	NAND_MUX_4x1 mux2_46(.out(stage3[46]), .select(sel[5:4]), .invSelect(invSel[5:4]), .in({{2{top}}, stage2[62], stage2[46]}));
	NAND_MUX_4x1 mux2_45(.out(stage3[45]), .select(sel[5:4]), .invSelect(invSel[5:4]), .in({{2{top}}, stage2[61], stage2[45]}));
	NAND_MUX_4x1 mux2_44(.out(stage3[44]), .select(sel[5:4]), .invSelect(invSel[5:4]), .in({{2{top}}, stage2[60], stage2[44]}));
	NAND_MUX_4x1 mux2_43(.out(stage3[43]), .select(sel[5:4]), .invSelect(invSel[5:4]), .in({{2{top}}, stage2[59], stage2[43]}));
	NAND_MUX_4x1 mux2_42(.out(stage3[42]), .select(sel[5:4]), .invSelect(invSel[5:4]), .in({{2{top}}, stage2[58], stage2[42]}));
	NAND_MUX_4x1 mux2_41(.out(stage3[41]), .select(sel[5:4]), .invSelect(invSel[5:4]), .in({{2{top}}, stage2[57], stage2[41]}));
	NAND_MUX_4x1 mux2_40(.out(stage3[40]), .select(sel[5:4]), .invSelect(invSel[5:4]), .in({{2{top}}, stage2[56], stage2[40]}));
		NAND_MUX_4x1 mux2_55(.out(stage3[55]), .select(sel[5:4]), .invSelect(invSel[5:4]), .in({{3{top}}, stage2[55]}));
	NAND_MUX_4x1 mux2_54(.out(stage3[54]), .select(sel[5:4]), .invSelect(invSel[5:4]), .in({{3{top}}, stage2[54]}));
	NAND_MUX_4x1 mux2_53(.out(stage3[53]), .select(sel[5:4]), .invSelect(invSel[5:4]), .in({{3{top}}, stage2[53]}));
	NAND_MUX_4x1 mux2_52(.out(stage3[52]), .select(sel[5:4]), .invSelect(invSel[5:4]), .in({{3{top}}, stage2[52]}));
	NAND_MUX_4x1 mux2_51(.out(stage3[51]), .select(sel[5:4]), .invSelect(invSel[5:4]), .in({{3{top}}, stage2[51]}));
	NAND_MUX_4x1 mux2_50(.out(stage3[50]), .select(sel[5:4]), .invSelect(invSel[5:4]), .in({{3{top}}, stage2[50]}));
	NAND_MUX_4x1 mux2_49(.out(stage3[49]), .select(sel[5:4]), .invSelect(invSel[5:4]), .in({{3{top}}, stage2[49]}));
	NAND_MUX_4x1 mux2_48(.out(stage3[48]), .select(sel[5:4]), .invSelect(invSel[5:4]), .in({{3{top}}, stage2[48]}));
		NAND_MUX_4x1 mux2_63(.out(stage3[63]), .select(sel[5:4]), .invSelect(invSel[5:4]), .in({{3{top}}, stage2[63]}));
	NAND_MUX_4x1 mux2_62(.out(stage3[62]), .select(sel[5:4]), .invSelect(invSel[5:4]), .in({{3{top}}, stage2[62]}));
	NAND_MUX_4x1 mux2_61(.out(stage3[61]), .select(sel[5:4]), .invSelect(invSel[5:4]), .in({{3{top}}, stage2[61]}));
	NAND_MUX_4x1 mux2_60(.out(stage3[60]), .select(sel[5:4]), .invSelect(invSel[5:4]), .in({{3{top}}, stage2[60]}));
	NAND_MUX_4x1 mux2_59(.out(stage3[59]), .select(sel[5:4]), .invSelect(invSel[5:4]), .in({{3{top}}, stage2[59]}));
	NAND_MUX_4x1 mux2_58(.out(stage3[58]), .select(sel[5:4]), .invSelect(invSel[5:4]), .in({{3{top}}, stage2[58]}));
	NAND_MUX_4x1 mux2_57(.out(stage3[57]), .select(sel[5:4]), .invSelect(invSel[5:4]), .in({{3{top}}, stage2[57]}));
	NAND_MUX_4x1 mux2_56(.out(stage3[56]), .select(sel[5:4]), .invSelect(invSel[5:4]), .in({{3{top}}, stage2[56]}));
	
	//stage 4, back to 63-0
		NAND_MUX_2x1 mux3_7(.out(out[7]), .select(left), .invSelect(invLeft), .in({stage3[-56], stage3[7]}));
	NAND_MUX_2x1 mux3_6(.out(out[6]), .select(left), .invSelect(invLeft), .in({stage3[-57], stage3[6]}));
	NAND_MUX_2x1 mux3_5(.out(out[5]), .select(left), .invSelect(invLeft), .in({stage3[-58], stage3[5]}));
	NAND_MUX_2x1 mux3_4(.out(out[4]), .select(left), .invSelect(invLeft), .in({stage3[-59], stage3[4]}));
	NAND_MUX_2x1 mux3_3(.out(out[3]), .select(left), .invSelect(invLeft), .in({stage3[-60], stage3[3]}));
	NAND_MUX_2x1 mux3_2(.out(out[2]), .select(left), .invSelect(invLeft), .in({stage3[-61], stage3[2]}));
	NAND_MUX_2x1 mux3_1(.out(out[1]), .select(left), .invSelect(invLeft), .in({stage3[-62], stage3[1]}));
	NAND_MUX_2x1 mux3_0(.out(out[0]), .select(left), .invSelect(invLeft), .in({stage3[-63], stage3[0]}));
		NAND_MUX_2x1 mux3_15(.out(out[15]), .select(left), .invSelect(invLeft), .in({stage3[-48], stage3[15]}));
	NAND_MUX_2x1 mux3_14(.out(out[14]), .select(left), .invSelect(invLeft), .in({stage3[-49], stage3[14]}));
	NAND_MUX_2x1 mux3_13(.out(out[13]), .select(left), .invSelect(invLeft), .in({stage3[-50], stage3[13]}));
	NAND_MUX_2x1 mux3_12(.out(out[12]), .select(left), .invSelect(invLeft), .in({stage3[-51], stage3[12]}));
	NAND_MUX_2x1 mux3_11(.out(out[11]), .select(left), .invSelect(invLeft), .in({stage3[-52], stage3[11]}));
	NAND_MUX_2x1 mux3_10(.out(out[10]), .select(left), .invSelect(invLeft), .in({stage3[-53], stage3[10]}));
	NAND_MUX_2x1 mux3_9(.out(out[9]), .select(left), .invSelect(invLeft), .in({stage3[-54], stage3[9]}));
	NAND_MUX_2x1 mux3_8(.out(out[8]), .select(left), .invSelect(invLeft), .in({stage3[-55], stage3[8]}));
		NAND_MUX_2x1 mux3_23(.out(out[23]), .select(left), .invSelect(invLeft), .in({stage3[-40], stage3[23]}));
	NAND_MUX_2x1 mux3_22(.out(out[22]), .select(left), .invSelect(invLeft), .in({stage3[-41], stage3[22]}));
	NAND_MUX_2x1 mux3_21(.out(out[21]), .select(left), .invSelect(invLeft), .in({stage3[-42], stage3[21]}));
	NAND_MUX_2x1 mux3_20(.out(out[20]), .select(left), .invSelect(invLeft), .in({stage3[-43], stage3[20]}));
	NAND_MUX_2x1 mux3_19(.out(out[19]), .select(left), .invSelect(invLeft), .in({stage3[-44], stage3[19]}));
	NAND_MUX_2x1 mux3_18(.out(out[18]), .select(left), .invSelect(invLeft), .in({stage3[-45], stage3[18]}));
	NAND_MUX_2x1 mux3_17(.out(out[17]), .select(left), .invSelect(invLeft), .in({stage3[-46], stage3[17]}));
	NAND_MUX_2x1 mux3_16(.out(out[16]), .select(left), .invSelect(invLeft), .in({stage3[-47], stage3[16]}));
		NAND_MUX_2x1 mux3_31(.out(out[31]), .select(left), .invSelect(invLeft), .in({stage3[-32], stage3[31]}));
	NAND_MUX_2x1 mux3_30(.out(out[30]), .select(left), .invSelect(invLeft), .in({stage3[-33], stage3[30]}));
	NAND_MUX_2x1 mux3_29(.out(out[29]), .select(left), .invSelect(invLeft), .in({stage3[-34], stage3[29]}));
	NAND_MUX_2x1 mux3_28(.out(out[28]), .select(left), .invSelect(invLeft), .in({stage3[-35], stage3[28]}));
	NAND_MUX_2x1 mux3_27(.out(out[27]), .select(left), .invSelect(invLeft), .in({stage3[-36], stage3[27]}));
	NAND_MUX_2x1 mux3_26(.out(out[26]), .select(left), .invSelect(invLeft), .in({stage3[-37], stage3[26]}));
	NAND_MUX_2x1 mux3_25(.out(out[25]), .select(left), .invSelect(invLeft), .in({stage3[-38], stage3[25]}));
	NAND_MUX_2x1 mux3_24(.out(out[24]), .select(left), .invSelect(invLeft), .in({stage3[-39], stage3[24]}));
		NAND_MUX_2x1 mux3_39(.out(out[39]), .select(left), .invSelect(invLeft), .in({stage3[-24], stage3[39]}));
	NAND_MUX_2x1 mux3_38(.out(out[38]), .select(left), .invSelect(invLeft), .in({stage3[-25], stage3[38]}));
	NAND_MUX_2x1 mux3_37(.out(out[37]), .select(left), .invSelect(invLeft), .in({stage3[-26], stage3[37]}));
	NAND_MUX_2x1 mux3_36(.out(out[36]), .select(left), .invSelect(invLeft), .in({stage3[-27], stage3[36]}));
	NAND_MUX_2x1 mux3_35(.out(out[35]), .select(left), .invSelect(invLeft), .in({stage3[-28], stage3[35]}));
	NAND_MUX_2x1 mux3_34(.out(out[34]), .select(left), .invSelect(invLeft), .in({stage3[-29], stage3[34]}));
	NAND_MUX_2x1 mux3_33(.out(out[33]), .select(left), .invSelect(invLeft), .in({stage3[-30], stage3[33]}));
	NAND_MUX_2x1 mux3_32(.out(out[32]), .select(left), .invSelect(invLeft), .in({stage3[-31], stage3[32]}));
		NAND_MUX_2x1 mux3_47(.out(out[47]), .select(left), .invSelect(invLeft), .in({stage3[-16], stage3[47]}));
	NAND_MUX_2x1 mux3_46(.out(out[46]), .select(left), .invSelect(invLeft), .in({stage3[-17], stage3[46]}));
	NAND_MUX_2x1 mux3_45(.out(out[45]), .select(left), .invSelect(invLeft), .in({stage3[-18], stage3[45]}));
	NAND_MUX_2x1 mux3_44(.out(out[44]), .select(left), .invSelect(invLeft), .in({stage3[-19], stage3[44]}));
	NAND_MUX_2x1 mux3_43(.out(out[43]), .select(left), .invSelect(invLeft), .in({stage3[-20], stage3[43]}));
	NAND_MUX_2x1 mux3_42(.out(out[42]), .select(left), .invSelect(invLeft), .in({stage3[-21], stage3[42]}));
	NAND_MUX_2x1 mux3_41(.out(out[41]), .select(left), .invSelect(invLeft), .in({stage3[-22], stage3[41]}));
	NAND_MUX_2x1 mux3_40(.out(out[40]), .select(left), .invSelect(invLeft), .in({stage3[-23], stage3[40]}));
		NAND_MUX_2x1 mux3_55(.out(out[55]), .select(left), .invSelect(invLeft), .in({stage3[-8], stage3[55]}));
	NAND_MUX_2x1 mux3_54(.out(out[54]), .select(left), .invSelect(invLeft), .in({stage3[-9], stage3[54]}));
	NAND_MUX_2x1 mux3_53(.out(out[53]), .select(left), .invSelect(invLeft), .in({stage3[-10], stage3[53]}));
	NAND_MUX_2x1 mux3_52(.out(out[52]), .select(left), .invSelect(invLeft), .in({stage3[-11], stage3[52]}));
	NAND_MUX_2x1 mux3_51(.out(out[51]), .select(left), .invSelect(invLeft), .in({stage3[-12], stage3[51]}));
	NAND_MUX_2x1 mux3_50(.out(out[50]), .select(left), .invSelect(invLeft), .in({stage3[-13], stage3[50]}));
	NAND_MUX_2x1 mux3_49(.out(out[49]), .select(left), .invSelect(invLeft), .in({stage3[-14], stage3[49]}));
	NAND_MUX_2x1 mux3_48(.out(out[48]), .select(left), .invSelect(invLeft), .in({stage3[-15], stage3[48]}));
		NAND_MUX_2x1 mux3_63(.out(out[63]), .select(left), .invSelect(invLeft), .in({stage3[0], stage3[63]}));
	NAND_MUX_2x1 mux3_62(.out(out[62]), .select(left), .invSelect(invLeft), .in({stage3[-1], stage3[62]}));
	NAND_MUX_2x1 mux3_61(.out(out[61]), .select(left), .invSelect(invLeft), .in({stage3[-2], stage3[61]}));
	NAND_MUX_2x1 mux3_60(.out(out[60]), .select(left), .invSelect(invLeft), .in({stage3[-3], stage3[60]}));
	NAND_MUX_2x1 mux3_59(.out(out[59]), .select(left), .invSelect(invLeft), .in({stage3[-4], stage3[59]}));
	NAND_MUX_2x1 mux3_58(.out(out[58]), .select(left), .invSelect(invLeft), .in({stage3[-5], stage3[58]}));
	NAND_MUX_2x1 mux3_57(.out(out[57]), .select(left), .invSelect(invLeft), .in({stage3[-6], stage3[57]}));
	NAND_MUX_2x1 mux3_56(.out(out[56]), .select(left), .invSelect(invLeft), .in({stage3[-7], stage3[56]}));
endmodule

/*
module shifter_testbench;
	wire [63:0] out;
	reg [5:0] shamt;
	reg left, sign;
	reg [63:0] in;
	shifter dut(.out, .shamt, .left, .sign, .in);
	assign sign=0; //no sign extend for now
	
	initial begin
	in = 64'h0000_0000_0000_0000;
	shamt = 6'h00;
	left=0;
	#10;
	in = 64'hF123_4567_89AB_CDEF;
	#10;
	shamt=6'h4;
	#10;
	shamt=6'h10;
	#10;
	shamt=6'h13;
	#10;
	shamt=6'h8;
	left=1;
	#10;
	shamt=6'h12;
	#10;
	shamt=6'h3F;
	#10;
	left=0;
	#10;
	end
endmodule */

