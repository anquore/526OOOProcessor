module fullAdderArray63(S, Cout, A, B, Cin);
	output [62:0] S, Cout;
	input [62:0] A, B, Cin;
	
		full_adder add7(.S(S[7]), .Cout(Cout[7]), .A(A[7]), .B(B[7]), .Cin(Cin[7]));
	full_adder add6(.S(S[6]), .Cout(Cout[6]), .A(A[6]), .B(B[6]), .Cin(Cin[6]));
	full_adder add5(.S(S[5]), .Cout(Cout[5]), .A(A[5]), .B(B[5]), .Cin(Cin[5]));
	full_adder add4(.S(S[4]), .Cout(Cout[4]), .A(A[4]), .B(B[4]), .Cin(Cin[4]));
	full_adder add3(.S(S[3]), .Cout(Cout[3]), .A(A[3]), .B(B[3]), .Cin(Cin[3]));
	full_adder add2(.S(S[2]), .Cout(Cout[2]), .A(A[2]), .B(B[2]), .Cin(Cin[2]));
	full_adder add1(.S(S[1]), .Cout(Cout[1]), .A(A[1]), .B(B[1]), .Cin(Cin[1]));
	full_adder add0(.S(S[0]), .Cout(Cout[0]), .A(A[0]), .B(B[0]), .Cin(Cin[0]));
		full_adder add15(.S(S[15]), .Cout(Cout[15]), .A(A[15]), .B(B[15]), .Cin(Cin[15]));
	full_adder add14(.S(S[14]), .Cout(Cout[14]), .A(A[14]), .B(B[14]), .Cin(Cin[14]));
	full_adder add13(.S(S[13]), .Cout(Cout[13]), .A(A[13]), .B(B[13]), .Cin(Cin[13]));
	full_adder add12(.S(S[12]), .Cout(Cout[12]), .A(A[12]), .B(B[12]), .Cin(Cin[12]));
	full_adder add11(.S(S[11]), .Cout(Cout[11]), .A(A[11]), .B(B[11]), .Cin(Cin[11]));
	full_adder add10(.S(S[10]), .Cout(Cout[10]), .A(A[10]), .B(B[10]), .Cin(Cin[10]));
	full_adder add9(.S(S[9]), .Cout(Cout[9]), .A(A[9]), .B(B[9]), .Cin(Cin[9]));
	full_adder add8(.S(S[8]), .Cout(Cout[8]), .A(A[8]), .B(B[8]), .Cin(Cin[8]));
		full_adder add23(.S(S[23]), .Cout(Cout[23]), .A(A[23]), .B(B[23]), .Cin(Cin[23]));
	full_adder add22(.S(S[22]), .Cout(Cout[22]), .A(A[22]), .B(B[22]), .Cin(Cin[22]));
	full_adder add21(.S(S[21]), .Cout(Cout[21]), .A(A[21]), .B(B[21]), .Cin(Cin[21]));
	full_adder add20(.S(S[20]), .Cout(Cout[20]), .A(A[20]), .B(B[20]), .Cin(Cin[20]));
	full_adder add19(.S(S[19]), .Cout(Cout[19]), .A(A[19]), .B(B[19]), .Cin(Cin[19]));
	full_adder add18(.S(S[18]), .Cout(Cout[18]), .A(A[18]), .B(B[18]), .Cin(Cin[18]));
	full_adder add17(.S(S[17]), .Cout(Cout[17]), .A(A[17]), .B(B[17]), .Cin(Cin[17]));
	full_adder add16(.S(S[16]), .Cout(Cout[16]), .A(A[16]), .B(B[16]), .Cin(Cin[16]));
		full_adder add31(.S(S[31]), .Cout(Cout[31]), .A(A[31]), .B(B[31]), .Cin(Cin[31]));
	full_adder add30(.S(S[30]), .Cout(Cout[30]), .A(A[30]), .B(B[30]), .Cin(Cin[30]));
	full_adder add29(.S(S[29]), .Cout(Cout[29]), .A(A[29]), .B(B[29]), .Cin(Cin[29]));
	full_adder add28(.S(S[28]), .Cout(Cout[28]), .A(A[28]), .B(B[28]), .Cin(Cin[28]));
	full_adder add27(.S(S[27]), .Cout(Cout[27]), .A(A[27]), .B(B[27]), .Cin(Cin[27]));
	full_adder add26(.S(S[26]), .Cout(Cout[26]), .A(A[26]), .B(B[26]), .Cin(Cin[26]));
	full_adder add25(.S(S[25]), .Cout(Cout[25]), .A(A[25]), .B(B[25]), .Cin(Cin[25]));
	full_adder add24(.S(S[24]), .Cout(Cout[24]), .A(A[24]), .B(B[24]), .Cin(Cin[24]));
		full_adder add39(.S(S[39]), .Cout(Cout[39]), .A(A[39]), .B(B[39]), .Cin(Cin[39]));
	full_adder add38(.S(S[38]), .Cout(Cout[38]), .A(A[38]), .B(B[38]), .Cin(Cin[38]));
	full_adder add37(.S(S[37]), .Cout(Cout[37]), .A(A[37]), .B(B[37]), .Cin(Cin[37]));
	full_adder add36(.S(S[36]), .Cout(Cout[36]), .A(A[36]), .B(B[36]), .Cin(Cin[36]));
	full_adder add35(.S(S[35]), .Cout(Cout[35]), .A(A[35]), .B(B[35]), .Cin(Cin[35]));
	full_adder add34(.S(S[34]), .Cout(Cout[34]), .A(A[34]), .B(B[34]), .Cin(Cin[34]));
	full_adder add33(.S(S[33]), .Cout(Cout[33]), .A(A[33]), .B(B[33]), .Cin(Cin[33]));
	full_adder add32(.S(S[32]), .Cout(Cout[32]), .A(A[32]), .B(B[32]), .Cin(Cin[32]));
		full_adder add47(.S(S[47]), .Cout(Cout[47]), .A(A[47]), .B(B[47]), .Cin(Cin[47]));
	full_adder add46(.S(S[46]), .Cout(Cout[46]), .A(A[46]), .B(B[46]), .Cin(Cin[46]));
	full_adder add45(.S(S[45]), .Cout(Cout[45]), .A(A[45]), .B(B[45]), .Cin(Cin[45]));
	full_adder add44(.S(S[44]), .Cout(Cout[44]), .A(A[44]), .B(B[44]), .Cin(Cin[44]));
	full_adder add43(.S(S[43]), .Cout(Cout[43]), .A(A[43]), .B(B[43]), .Cin(Cin[43]));
	full_adder add42(.S(S[42]), .Cout(Cout[42]), .A(A[42]), .B(B[42]), .Cin(Cin[42]));
	full_adder add41(.S(S[41]), .Cout(Cout[41]), .A(A[41]), .B(B[41]), .Cin(Cin[41]));
	full_adder add40(.S(S[40]), .Cout(Cout[40]), .A(A[40]), .B(B[40]), .Cin(Cin[40]));
		full_adder add55(.S(S[55]), .Cout(Cout[55]), .A(A[55]), .B(B[55]), .Cin(Cin[55]));
	full_adder add54(.S(S[54]), .Cout(Cout[54]), .A(A[54]), .B(B[54]), .Cin(Cin[54]));
	full_adder add53(.S(S[53]), .Cout(Cout[53]), .A(A[53]), .B(B[53]), .Cin(Cin[53]));
	full_adder add52(.S(S[52]), .Cout(Cout[52]), .A(A[52]), .B(B[52]), .Cin(Cin[52]));
	full_adder add51(.S(S[51]), .Cout(Cout[51]), .A(A[51]), .B(B[51]), .Cin(Cin[51]));
	full_adder add50(.S(S[50]), .Cout(Cout[50]), .A(A[50]), .B(B[50]), .Cin(Cin[50]));
	full_adder add49(.S(S[49]), .Cout(Cout[49]), .A(A[49]), .B(B[49]), .Cin(Cin[49]));
	full_adder add48(.S(S[48]), .Cout(Cout[48]), .A(A[48]), .B(B[48]), .Cin(Cin[48]));
	
	full_adder add62(.S(S[62]), .Cout(Cout[62]), .A(A[62]), .B(B[62]), .Cin(Cin[62]));
	full_adder add61(.S(S[61]), .Cout(Cout[61]), .A(A[61]), .B(B[61]), .Cin(Cin[51]));
	full_adder add60(.S(S[60]), .Cout(Cout[60]), .A(A[60]), .B(B[60]), .Cin(Cin[60]));
	full_adder add59(.S(S[59]), .Cout(Cout[59]), .A(A[59]), .B(B[59]), .Cin(Cin[59]));
	full_adder add58(.S(S[58]), .Cout(Cout[58]), .A(A[58]), .B(B[58]), .Cin(Cin[58]));
	full_adder add57(.S(S[57]), .Cout(Cout[57]), .A(A[57]), .B(B[57]), .Cin(Cin[57]));
	full_adder add56(.S(S[56]), .Cout(Cout[56]), .A(A[56]), .B(B[56]), .Cin(Cin[56]));
endmodule
