module mux16x1X64(outs, addr, muxIns);
	output [63:0] outs;
	input [3:0] addr;
	input [15:0][63:0] muxIns;
	
	mux16x1 mux7(.out(outs[7]), .addr, .muxIns({muxIns[15][7], muxIns[14][7], muxIns[13][7], muxIns[12][7], muxIns[11][7], muxIns[10][7], muxIns[9][7], muxIns[8][7],
		muxIns[7][7], muxIns[6][7], muxIns[5][7], muxIns[4][7], muxIns[3][7], muxIns[2][7], muxIns[1][7], muxIns[0][7]}));
	mux16x1 mux6(.out(outs[6]), .addr, .muxIns({muxIns[15][6], muxIns[14][6], muxIns[13][6], muxIns[12][6], muxIns[11][6], muxIns[10][6], muxIns[9][6], muxIns[8][6],
		muxIns[7][6], muxIns[6][6], muxIns[5][6], muxIns[4][6], muxIns[3][6], muxIns[2][6], muxIns[1][6], muxIns[0][6]}));
	mux16x1 mux5(.out(outs[5]), .addr, .muxIns({muxIns[15][5], muxIns[14][5], muxIns[13][5], muxIns[12][5], muxIns[11][5], muxIns[10][5], muxIns[9][5], muxIns[8][5],
		muxIns[7][5], muxIns[6][5], muxIns[5][5], muxIns[4][5], muxIns[3][5], muxIns[2][5], muxIns[1][5], muxIns[0][5]}));
	mux16x1 mux4(.out(outs[4]), .addr, .muxIns({muxIns[15][4], muxIns[14][4], muxIns[13][4], muxIns[12][4], muxIns[11][4], muxIns[10][4], muxIns[9][4], muxIns[8][4],
		muxIns[7][4], muxIns[6][4], muxIns[5][4], muxIns[4][4], muxIns[3][4], muxIns[2][4], muxIns[1][4], muxIns[0][4]}));
	mux16x1 mux3(.out(outs[3]), .addr, .muxIns({muxIns[15][3], muxIns[14][3], muxIns[13][3], muxIns[12][3], muxIns[11][3], muxIns[10][3], muxIns[9][3], muxIns[8][3],
		muxIns[7][3], muxIns[6][3], muxIns[5][3], muxIns[4][3], muxIns[3][3], muxIns[2][3], muxIns[1][3], muxIns[0][3]}));
	mux16x1 mux2(.out(outs[2]), .addr, .muxIns({muxIns[15][2], muxIns[14][2], muxIns[13][2], muxIns[12][2], muxIns[11][2], muxIns[10][2], muxIns[9][2], muxIns[8][2],
		muxIns[7][2], muxIns[6][2], muxIns[5][2], muxIns[4][2], muxIns[3][2], muxIns[2][2], muxIns[1][2], muxIns[0][2]}));
	mux16x1 mux1(.out(outs[1]), .addr, .muxIns({muxIns[15][1], muxIns[14][1], muxIns[13][1], muxIns[12][1], muxIns[11][1], muxIns[10][1], muxIns[9][1], muxIns[8][1],
		muxIns[7][1], muxIns[6][1], muxIns[5][1], muxIns[4][1], muxIns[3][1], muxIns[2][1], muxIns[1][1], muxIns[0][1]}));
	mux16x1 mux0(.out(outs[0]), .addr, .muxIns({muxIns[15][0], muxIns[14][0], muxIns[13][0], muxIns[12][0], muxIns[11][0], muxIns[10][0], muxIns[9][0], muxIns[8][0],
		muxIns[7][0], muxIns[6][0], muxIns[5][0], muxIns[4][0], muxIns[3][0], muxIns[2][0], muxIns[1][0], muxIns[0][0]}));
	
	mux16x1 mux15(.out(outs[15]), .addr, .muxIns({muxIns[15][15], muxIns[14][15], muxIns[13][15], muxIns[12][15], muxIns[11][15], muxIns[10][15], muxIns[9][15], muxIns[8][15],
		muxIns[7][15], muxIns[6][15], muxIns[5][15], muxIns[4][15], muxIns[3][15], muxIns[2][15], muxIns[1][15], muxIns[0][15]}));
	mux16x1 mux14(.out(outs[14]), .addr, .muxIns({muxIns[15][14], muxIns[14][14], muxIns[13][14], muxIns[12][14], muxIns[11][14], muxIns[10][14], muxIns[9][14], muxIns[8][14],
		muxIns[7][14], muxIns[6][14], muxIns[5][14], muxIns[4][14], muxIns[3][14], muxIns[2][14], muxIns[1][14], muxIns[0][14]}));
	mux16x1 mux13(.out(outs[13]), .addr, .muxIns({muxIns[15][13], muxIns[14][13], muxIns[13][13], muxIns[12][13], muxIns[11][13], muxIns[10][13], muxIns[9][13], muxIns[8][13],
		muxIns[7][13], muxIns[6][13], muxIns[5][13], muxIns[4][13], muxIns[3][13], muxIns[2][13], muxIns[1][13], muxIns[0][13]}));
	mux16x1 mux12(.out(outs[12]), .addr, .muxIns({muxIns[15][12], muxIns[14][12], muxIns[13][12], muxIns[12][12], muxIns[11][12], muxIns[10][12], muxIns[9][12], muxIns[8][12],
		muxIns[7][12], muxIns[6][12], muxIns[5][12], muxIns[4][12], muxIns[3][12], muxIns[2][12], muxIns[1][12], muxIns[0][12]}));
	mux16x1 mux11(.out(outs[11]), .addr, .muxIns({muxIns[15][11], muxIns[14][11], muxIns[13][11], muxIns[12][11], muxIns[11][11], muxIns[10][11], muxIns[9][11], muxIns[8][11],
		muxIns[7][11], muxIns[6][11], muxIns[5][11], muxIns[4][11], muxIns[3][11], muxIns[2][11], muxIns[1][11], muxIns[0][11]}));
	mux16x1 mux10(.out(outs[10]), .addr, .muxIns({muxIns[15][10], muxIns[14][10], muxIns[13][10], muxIns[12][10], muxIns[11][10], muxIns[10][10], muxIns[9][10], muxIns[8][10],
		muxIns[7][10], muxIns[6][10], muxIns[5][10], muxIns[4][10], muxIns[3][10], muxIns[2][10], muxIns[1][10], muxIns[0][10]}));
	mux16x1 mux9(.out(outs[9]), .addr, .muxIns({muxIns[15][9], muxIns[14][9], muxIns[13][9], muxIns[12][9], muxIns[11][9], muxIns[10][9], muxIns[9][9], muxIns[8][9],
		muxIns[7][9], muxIns[6][9], muxIns[5][9], muxIns[4][9], muxIns[3][9], muxIns[2][9], muxIns[1][9], muxIns[0][9]}));
	mux16x1 mux8(.out(outs[8]), .addr, .muxIns({muxIns[15][8], muxIns[14][8], muxIns[13][8], muxIns[12][8], muxIns[11][8], muxIns[10][8], muxIns[9][8], muxIns[8][8],
		muxIns[7][8], muxIns[6][8], muxIns[5][8], muxIns[4][8], muxIns[3][8], muxIns[2][8], muxIns[1][8], muxIns[0][8]}));
	
	mux16x1 mux23(.out(outs[23]), .addr, .muxIns({muxIns[15][23], muxIns[14][23], muxIns[13][23], muxIns[12][23], muxIns[11][23], muxIns[10][23], muxIns[9][23], muxIns[8][23],
		muxIns[7][23], muxIns[6][23], muxIns[5][23], muxIns[4][23], muxIns[3][23], muxIns[2][23], muxIns[1][23], muxIns[0][23]}));
	mux16x1 mux22(.out(outs[22]), .addr, .muxIns({muxIns[15][22], muxIns[14][22], muxIns[13][22], muxIns[12][22], muxIns[11][22], muxIns[10][22], muxIns[9][22], muxIns[8][22],
		muxIns[7][22], muxIns[6][22], muxIns[5][22], muxIns[4][22], muxIns[3][22], muxIns[2][22], muxIns[1][22], muxIns[0][22]}));
	mux16x1 mux21(.out(outs[21]), .addr, .muxIns({muxIns[15][21], muxIns[14][21], muxIns[13][21], muxIns[12][21], muxIns[11][21], muxIns[10][21], muxIns[9][21], muxIns[8][21],
		muxIns[7][21], muxIns[6][21], muxIns[5][21], muxIns[4][21], muxIns[3][21], muxIns[2][21], muxIns[1][21], muxIns[0][21]}));
	mux16x1 mux20(.out(outs[20]), .addr, .muxIns({muxIns[15][20], muxIns[14][20], muxIns[13][20], muxIns[12][20], muxIns[11][20], muxIns[10][20], muxIns[9][20], muxIns[8][20],
		muxIns[7][20], muxIns[6][20], muxIns[5][20], muxIns[4][20], muxIns[3][20], muxIns[2][20], muxIns[1][20], muxIns[0][20]}));
	mux16x1 mux19(.out(outs[19]), .addr, .muxIns({muxIns[15][19], muxIns[14][19], muxIns[13][19], muxIns[12][19], muxIns[11][19], muxIns[10][19], muxIns[9][19], muxIns[8][19],
		muxIns[7][19], muxIns[6][19], muxIns[5][19], muxIns[4][19], muxIns[3][19], muxIns[2][19], muxIns[1][19], muxIns[0][19]}));
	mux16x1 mux18(.out(outs[18]), .addr, .muxIns({muxIns[15][18], muxIns[14][18], muxIns[13][18], muxIns[12][18], muxIns[11][18], muxIns[10][18], muxIns[9][18], muxIns[8][18],
		muxIns[7][18], muxIns[6][18], muxIns[5][18], muxIns[4][18], muxIns[3][18], muxIns[2][18], muxIns[1][18], muxIns[0][18]}));
	mux16x1 mux17(.out(outs[17]), .addr, .muxIns({muxIns[15][17], muxIns[14][17], muxIns[13][17], muxIns[12][17], muxIns[11][17], muxIns[10][17], muxIns[9][17], muxIns[8][17],
		muxIns[7][17], muxIns[6][17], muxIns[5][17], muxIns[4][17], muxIns[3][17], muxIns[2][17], muxIns[1][17], muxIns[0][17]}));
	mux16x1 mux16(.out(outs[16]), .addr, .muxIns({muxIns[15][16], muxIns[14][16], muxIns[13][16], muxIns[12][16], muxIns[11][16], muxIns[10][16], muxIns[9][16], muxIns[8][16],
		muxIns[7][16], muxIns[6][16], muxIns[5][16], muxIns[4][16], muxIns[3][16], muxIns[2][16], muxIns[1][16], muxIns[0][16]}));
	
	mux16x1 mux31(.out(outs[31]), .addr, .muxIns({muxIns[15][31], muxIns[14][31], muxIns[13][31], muxIns[12][31], muxIns[11][31], muxIns[10][31], muxIns[9][31], muxIns[8][31],
		muxIns[7][31], muxIns[6][31], muxIns[5][31], muxIns[4][31], muxIns[3][31], muxIns[2][31], muxIns[1][31], muxIns[0][31]}));
	mux16x1 mux30(.out(outs[30]), .addr, .muxIns({muxIns[15][30], muxIns[14][30], muxIns[13][30], muxIns[12][30], muxIns[11][30], muxIns[10][30], muxIns[9][30], muxIns[8][30],
		muxIns[7][30], muxIns[6][30], muxIns[5][30], muxIns[4][30], muxIns[3][30], muxIns[2][30], muxIns[1][30], muxIns[0][30]}));
	mux16x1 mux29(.out(outs[29]), .addr, .muxIns({muxIns[15][29], muxIns[14][29], muxIns[13][29], muxIns[12][29], muxIns[11][29], muxIns[10][29], muxIns[9][29], muxIns[8][29],
		muxIns[7][29], muxIns[6][29], muxIns[5][29], muxIns[4][29], muxIns[3][29], muxIns[2][29], muxIns[1][29], muxIns[0][29]}));
	mux16x1 mux28(.out(outs[28]), .addr, .muxIns({muxIns[15][28], muxIns[14][28], muxIns[13][28], muxIns[12][28], muxIns[11][28], muxIns[10][28], muxIns[9][28], muxIns[8][28],
		muxIns[7][28], muxIns[6][28], muxIns[5][28], muxIns[4][28], muxIns[3][28], muxIns[2][28], muxIns[1][28], muxIns[0][28]}));
	mux16x1 mux27(.out(outs[27]), .addr, .muxIns({muxIns[15][27], muxIns[14][27], muxIns[13][27], muxIns[12][27], muxIns[11][27], muxIns[10][27], muxIns[9][27], muxIns[8][27],
		muxIns[7][27], muxIns[6][27], muxIns[5][27], muxIns[4][27], muxIns[3][27], muxIns[2][27], muxIns[1][27], muxIns[0][27]}));
	mux16x1 mux26(.out(outs[26]), .addr, .muxIns({muxIns[15][26], muxIns[14][26], muxIns[13][26], muxIns[12][26], muxIns[11][26], muxIns[10][26], muxIns[9][26], muxIns[8][26],
		muxIns[7][26], muxIns[6][26], muxIns[5][26], muxIns[4][26], muxIns[3][26], muxIns[2][26], muxIns[1][26], muxIns[0][26]}));
	mux16x1 mux25(.out(outs[25]), .addr, .muxIns({muxIns[15][25], muxIns[14][25], muxIns[13][25], muxIns[12][25], muxIns[11][25], muxIns[10][25], muxIns[9][25], muxIns[8][25],
		muxIns[7][25], muxIns[6][25], muxIns[5][25], muxIns[4][25], muxIns[3][25], muxIns[2][25], muxIns[1][25], muxIns[0][25]}));
	mux16x1 mux24(.out(outs[24]), .addr, .muxIns({muxIns[15][24], muxIns[14][24], muxIns[13][24], muxIns[12][24], muxIns[11][24], muxIns[10][24], muxIns[9][24], muxIns[8][24],
		muxIns[7][24], muxIns[6][24], muxIns[5][24], muxIns[4][24], muxIns[3][24], muxIns[2][24], muxIns[1][24], muxIns[0][24]}));
	
	mux16x1 mux39(.out(outs[39]), .addr, .muxIns({muxIns[15][39], muxIns[14][39], muxIns[13][39], muxIns[12][39], muxIns[11][39], muxIns[10][39], muxIns[9][39], muxIns[8][39],
		muxIns[7][39], muxIns[6][39], muxIns[5][39], muxIns[4][39], muxIns[3][39], muxIns[2][39], muxIns[1][39], muxIns[0][39]}));
	mux16x1 mux38(.out(outs[38]), .addr, .muxIns({muxIns[15][38], muxIns[14][38], muxIns[13][38], muxIns[12][38], muxIns[11][38], muxIns[10][38], muxIns[9][38], muxIns[8][38],
		muxIns[7][38], muxIns[6][38], muxIns[5][38], muxIns[4][38], muxIns[3][38], muxIns[2][38], muxIns[1][38], muxIns[0][38]}));
	mux16x1 mux37(.out(outs[37]), .addr, .muxIns({muxIns[15][37], muxIns[14][37], muxIns[13][37], muxIns[12][37], muxIns[11][37], muxIns[10][37], muxIns[9][37], muxIns[8][37],
		muxIns[7][37], muxIns[6][37], muxIns[5][37], muxIns[4][37], muxIns[3][37], muxIns[2][37], muxIns[1][37], muxIns[0][37]}));
	mux16x1 mux36(.out(outs[36]), .addr, .muxIns({muxIns[15][36], muxIns[14][36], muxIns[13][36], muxIns[12][36], muxIns[11][36], muxIns[10][36], muxIns[9][36], muxIns[8][36],
		muxIns[7][36], muxIns[6][36], muxIns[5][36], muxIns[4][36], muxIns[3][36], muxIns[2][36], muxIns[1][36], muxIns[0][36]}));
	mux16x1 mux35(.out(outs[35]), .addr, .muxIns({muxIns[15][35], muxIns[14][35], muxIns[13][35], muxIns[12][35], muxIns[11][35], muxIns[10][35], muxIns[9][35], muxIns[8][35],
		muxIns[7][35], muxIns[6][35], muxIns[5][35], muxIns[4][35], muxIns[3][35], muxIns[2][35], muxIns[1][35], muxIns[0][35]}));
	mux16x1 mux34(.out(outs[34]), .addr, .muxIns({muxIns[15][34], muxIns[14][34], muxIns[13][34], muxIns[12][34], muxIns[11][34], muxIns[10][34], muxIns[9][34], muxIns[8][34],
		muxIns[7][34], muxIns[6][34], muxIns[5][34], muxIns[4][34], muxIns[3][34], muxIns[2][34], muxIns[1][34], muxIns[0][34]}));
	mux16x1 mux33(.out(outs[33]), .addr, .muxIns({muxIns[15][33], muxIns[14][33], muxIns[13][33], muxIns[12][33], muxIns[11][33], muxIns[10][33], muxIns[9][33], muxIns[8][33],
		muxIns[7][33], muxIns[6][33], muxIns[5][33], muxIns[4][33], muxIns[3][33], muxIns[2][33], muxIns[1][33], muxIns[0][33]}));
	mux16x1 mux32(.out(outs[32]), .addr, .muxIns({muxIns[15][32], muxIns[14][32], muxIns[13][32], muxIns[12][32], muxIns[11][32], muxIns[10][32], muxIns[9][32], muxIns[8][32],
		muxIns[7][32], muxIns[6][32], muxIns[5][32], muxIns[4][32], muxIns[3][32], muxIns[2][32], muxIns[1][32], muxIns[0][32]}));
	
	mux16x1 mux47(.out(outs[47]), .addr, .muxIns({muxIns[15][47], muxIns[14][47], muxIns[13][47], muxIns[12][47], muxIns[11][47], muxIns[10][47], muxIns[9][47], muxIns[8][47],
		muxIns[7][47], muxIns[6][47], muxIns[5][47], muxIns[4][47], muxIns[3][47], muxIns[2][47], muxIns[1][47], muxIns[0][47]}));
	mux16x1 mux46(.out(outs[46]), .addr, .muxIns({muxIns[15][46], muxIns[14][46], muxIns[13][46], muxIns[12][46], muxIns[11][46], muxIns[10][46], muxIns[9][46], muxIns[8][46],
		muxIns[7][46], muxIns[6][46], muxIns[5][46], muxIns[4][46], muxIns[3][46], muxIns[2][46], muxIns[1][46], muxIns[0][46]}));
	mux16x1 mux45(.out(outs[45]), .addr, .muxIns({muxIns[15][45], muxIns[14][45], muxIns[13][45], muxIns[12][45], muxIns[11][45], muxIns[10][45], muxIns[9][45], muxIns[8][45],
		muxIns[7][45], muxIns[6][45], muxIns[5][45], muxIns[4][45], muxIns[3][45], muxIns[2][45], muxIns[1][45], muxIns[0][45]}));
	mux16x1 mux44(.out(outs[44]), .addr, .muxIns({muxIns[15][44], muxIns[14][44], muxIns[13][44], muxIns[12][44], muxIns[11][44], muxIns[10][44], muxIns[9][44], muxIns[8][44],
		muxIns[7][44], muxIns[6][44], muxIns[5][44], muxIns[4][44], muxIns[3][44], muxIns[2][44], muxIns[1][44], muxIns[0][44]}));
	mux16x1 mux43(.out(outs[43]), .addr, .muxIns({muxIns[15][43], muxIns[14][43], muxIns[13][43], muxIns[12][43], muxIns[11][43], muxIns[10][43], muxIns[9][43], muxIns[8][43],
		muxIns[7][43], muxIns[6][43], muxIns[5][43], muxIns[4][43], muxIns[3][43], muxIns[2][43], muxIns[1][43], muxIns[0][43]}));
	mux16x1 mux42(.out(outs[42]), .addr, .muxIns({muxIns[15][42], muxIns[14][42], muxIns[13][42], muxIns[12][42], muxIns[11][42], muxIns[10][42], muxIns[9][42], muxIns[8][42],
		muxIns[7][42], muxIns[6][42], muxIns[5][42], muxIns[4][42], muxIns[3][42], muxIns[2][42], muxIns[1][42], muxIns[0][42]}));
	mux16x1 mux41(.out(outs[41]), .addr, .muxIns({muxIns[15][41], muxIns[14][41], muxIns[13][41], muxIns[12][41], muxIns[11][41], muxIns[10][41], muxIns[9][41], muxIns[8][41],
		muxIns[7][41], muxIns[6][41], muxIns[5][41], muxIns[4][41], muxIns[3][41], muxIns[2][41], muxIns[1][41], muxIns[0][41]}));
	mux16x1 mux40(.out(outs[40]), .addr, .muxIns({muxIns[15][40], muxIns[14][40], muxIns[13][40], muxIns[12][40], muxIns[11][40], muxIns[10][40], muxIns[9][40], muxIns[8][40],
		muxIns[7][40], muxIns[6][40], muxIns[5][40], muxIns[4][40], muxIns[3][40], muxIns[2][40], muxIns[1][40], muxIns[0][40]}));
	
	mux16x1 mux55(.out(outs[55]), .addr, .muxIns({muxIns[15][55], muxIns[14][55], muxIns[13][55], muxIns[12][55], muxIns[11][55], muxIns[10][55], muxIns[9][55], muxIns[8][55],
		muxIns[7][55], muxIns[6][55], muxIns[5][55], muxIns[4][55], muxIns[3][55], muxIns[2][55], muxIns[1][55], muxIns[0][55]}));
	mux16x1 mux54(.out(outs[54]), .addr, .muxIns({muxIns[15][54], muxIns[14][54], muxIns[13][54], muxIns[12][54], muxIns[11][54], muxIns[10][54], muxIns[9][54], muxIns[8][54],
		muxIns[7][54], muxIns[6][54], muxIns[5][54], muxIns[4][54], muxIns[3][54], muxIns[2][54], muxIns[1][54], muxIns[0][54]}));
	mux16x1 mux53(.out(outs[53]), .addr, .muxIns({muxIns[15][53], muxIns[14][53], muxIns[13][53], muxIns[12][53], muxIns[11][53], muxIns[10][53], muxIns[9][53], muxIns[8][53],
		muxIns[7][53], muxIns[6][53], muxIns[5][53], muxIns[4][53], muxIns[3][53], muxIns[2][53], muxIns[1][53], muxIns[0][53]}));
	mux16x1 mux52(.out(outs[52]), .addr, .muxIns({muxIns[15][52], muxIns[14][52], muxIns[13][52], muxIns[12][52], muxIns[11][52], muxIns[10][52], muxIns[9][52], muxIns[8][52],
		muxIns[7][52], muxIns[6][52], muxIns[5][52], muxIns[4][52], muxIns[3][52], muxIns[2][52], muxIns[1][52], muxIns[0][52]}));
	mux16x1 mux51(.out(outs[51]), .addr, .muxIns({muxIns[15][51], muxIns[14][51], muxIns[13][51], muxIns[12][51], muxIns[11][51], muxIns[10][51], muxIns[9][51], muxIns[8][51],
		muxIns[7][51], muxIns[6][51], muxIns[5][51], muxIns[4][51], muxIns[3][51], muxIns[2][51], muxIns[1][51], muxIns[0][51]}));
	mux16x1 mux50(.out(outs[50]), .addr, .muxIns({muxIns[15][50], muxIns[14][50], muxIns[13][50], muxIns[12][50], muxIns[11][50], muxIns[10][50], muxIns[9][50], muxIns[8][50],
		muxIns[7][50], muxIns[6][50], muxIns[5][50], muxIns[4][50], muxIns[3][50], muxIns[2][50], muxIns[1][50], muxIns[0][50]}));
	mux16x1 mux49(.out(outs[49]), .addr, .muxIns({muxIns[15][49], muxIns[14][49], muxIns[13][49], muxIns[12][49], muxIns[11][49], muxIns[10][49], muxIns[9][49], muxIns[8][49],
		muxIns[7][49], muxIns[6][49], muxIns[5][49], muxIns[4][49], muxIns[3][49], muxIns[2][49], muxIns[1][49], muxIns[0][49]}));
	mux16x1 mux48(.out(outs[48]), .addr, .muxIns({muxIns[15][48], muxIns[14][48], muxIns[13][48], muxIns[12][48], muxIns[11][48], muxIns[10][48], muxIns[9][48], muxIns[8][48],
		muxIns[7][48], muxIns[6][48], muxIns[5][48], muxIns[4][48], muxIns[3][48], muxIns[2][48], muxIns[1][48], muxIns[0][48]}));
	
	mux16x1 mux63(.out(outs[63]), .addr, .muxIns({muxIns[15][63], muxIns[14][63], muxIns[13][63], muxIns[12][63], muxIns[11][63], muxIns[10][63], muxIns[9][63], muxIns[8][63],
		muxIns[7][63], muxIns[6][63], muxIns[5][63], muxIns[4][63], muxIns[3][63], muxIns[2][63], muxIns[1][63], muxIns[0][63]}));
	mux16x1 mux62(.out(outs[62]), .addr, .muxIns({muxIns[15][62], muxIns[14][62], muxIns[13][62], muxIns[12][62], muxIns[11][62], muxIns[10][62], muxIns[9][62], muxIns[8][62],
		muxIns[7][62], muxIns[6][62], muxIns[5][62], muxIns[4][62], muxIns[3][62], muxIns[2][62], muxIns[1][62], muxIns[0][62]}));
	mux16x1 mux61(.out(outs[61]), .addr, .muxIns({muxIns[15][61], muxIns[14][61], muxIns[13][61], muxIns[12][61], muxIns[11][61], muxIns[10][61], muxIns[9][61], muxIns[8][61],
		muxIns[7][61], muxIns[6][61], muxIns[5][61], muxIns[4][61], muxIns[3][61], muxIns[2][61], muxIns[1][61], muxIns[0][61]}));
	mux16x1 mux60(.out(outs[60]), .addr, .muxIns({muxIns[15][60], muxIns[14][60], muxIns[13][60], muxIns[12][60], muxIns[11][60], muxIns[10][60], muxIns[9][60], muxIns[8][60],
		muxIns[7][60], muxIns[6][60], muxIns[5][60], muxIns[4][60], muxIns[3][60], muxIns[2][60], muxIns[1][60], muxIns[0][60]}));
	mux16x1 mux59(.out(outs[59]), .addr, .muxIns({muxIns[15][59], muxIns[14][59], muxIns[13][59], muxIns[12][59], muxIns[11][59], muxIns[10][59], muxIns[9][59], muxIns[8][59],
		muxIns[7][59], muxIns[6][59], muxIns[5][59], muxIns[4][59], muxIns[3][59], muxIns[2][59], muxIns[1][59], muxIns[0][59]}));
	mux16x1 mux58(.out(outs[58]), .addr, .muxIns({muxIns[15][58], muxIns[14][58], muxIns[13][58], muxIns[12][58], muxIns[11][58], muxIns[10][58], muxIns[9][58], muxIns[8][58],
		muxIns[7][58], muxIns[6][58], muxIns[5][58], muxIns[4][58], muxIns[3][58], muxIns[2][58], muxIns[1][58], muxIns[0][58]}));
	mux16x1 mux57(.out(outs[57]), .addr, .muxIns({muxIns[15][57], muxIns[14][57], muxIns[13][57], muxIns[12][57], muxIns[11][57], muxIns[10][57], muxIns[9][57], muxIns[8][57],
		muxIns[7][57], muxIns[6][57], muxIns[5][57], muxIns[4][57], muxIns[3][57], muxIns[2][57], muxIns[1][57], muxIns[0][57]}));
	mux16x1 mux56(.out(outs[56]), .addr, .muxIns({muxIns[15][56], muxIns[14][56], muxIns[13][56], muxIns[12][56], muxIns[11][56], muxIns[10][56], muxIns[9][56], muxIns[8][56],
		muxIns[7][56], muxIns[6][56], muxIns[5][56], muxIns[4][56], muxIns[3][56], muxIns[2][56], muxIns[1][56], muxIns[0][56]}));
endmodule

