module registerX64(outs, ins, en, rst, clk);
	output [63:0] outs;
	input [63:0] ins;
	input en, rst, clk;
	
	
		FF_en r7(.q(outs[7]), .d(ins[7]), .en, .reset(rst), .clk);
	FF_en r6(.q(outs[6]), .d(ins[6]), .en, .reset(rst), .clk);
	FF_en r5(.q(outs[5]), .d(ins[5]), .en, .reset(rst), .clk);
	FF_en r4(.q(outs[4]), .d(ins[4]), .en, .reset(rst), .clk);
	FF_en r3(.q(outs[3]), .d(ins[3]), .en, .reset(rst), .clk);
	FF_en r2(.q(outs[2]), .d(ins[2]), .en, .reset(rst), .clk);
	FF_en r1(.q(outs[1]), .d(ins[1]), .en, .reset(rst), .clk);
	FF_en r0(.q(outs[0]), .d(ins[0]), .en, .reset(rst), .clk);
		FF_en r15(.q(outs[15]), .d(ins[15]), .en, .reset(rst), .clk);
	FF_en r14(.q(outs[14]), .d(ins[14]), .en, .reset(rst), .clk);
	FF_en r13(.q(outs[13]), .d(ins[13]), .en, .reset(rst), .clk);
	FF_en r12(.q(outs[12]), .d(ins[12]), .en, .reset(rst), .clk);
	FF_en r11(.q(outs[11]), .d(ins[11]), .en, .reset(rst), .clk);
	FF_en r10(.q(outs[10]), .d(ins[10]), .en, .reset(rst), .clk);
	FF_en r9(.q(outs[9]), .d(ins[9]), .en, .reset(rst), .clk);
	FF_en r8(.q(outs[8]), .d(ins[8]), .en, .reset(rst), .clk);
		FF_en r23(.q(outs[23]), .d(ins[23]), .en, .reset(rst), .clk);
	FF_en r22(.q(outs[22]), .d(ins[22]), .en, .reset(rst), .clk);
	FF_en r21(.q(outs[21]), .d(ins[21]), .en, .reset(rst), .clk);
	FF_en r20(.q(outs[20]), .d(ins[20]), .en, .reset(rst), .clk);
	FF_en r19(.q(outs[19]), .d(ins[19]), .en, .reset(rst), .clk);
	FF_en r18(.q(outs[18]), .d(ins[18]), .en, .reset(rst), .clk);
	FF_en r17(.q(outs[17]), .d(ins[17]), .en, .reset(rst), .clk);
	FF_en r16(.q(outs[16]), .d(ins[16]), .en, .reset(rst), .clk);
		FF_en r31(.q(outs[31]), .d(ins[31]), .en, .reset(rst), .clk);
	FF_en r30(.q(outs[30]), .d(ins[30]), .en, .reset(rst), .clk);
	FF_en r29(.q(outs[29]), .d(ins[29]), .en, .reset(rst), .clk);
	FF_en r28(.q(outs[28]), .d(ins[28]), .en, .reset(rst), .clk);
	FF_en r27(.q(outs[27]), .d(ins[27]), .en, .reset(rst), .clk);
	FF_en r26(.q(outs[26]), .d(ins[26]), .en, .reset(rst), .clk);
	FF_en r25(.q(outs[25]), .d(ins[25]), .en, .reset(rst), .clk);
	FF_en r24(.q(outs[24]), .d(ins[24]), .en, .reset(rst), .clk);
		FF_en r39(.q(outs[39]), .d(ins[39]), .en, .reset(rst), .clk);
	FF_en r38(.q(outs[38]), .d(ins[38]), .en, .reset(rst), .clk);
	FF_en r37(.q(outs[37]), .d(ins[37]), .en, .reset(rst), .clk);
	FF_en r36(.q(outs[36]), .d(ins[36]), .en, .reset(rst), .clk);
	FF_en r35(.q(outs[35]), .d(ins[35]), .en, .reset(rst), .clk);
	FF_en r34(.q(outs[34]), .d(ins[34]), .en, .reset(rst), .clk);
	FF_en r33(.q(outs[33]), .d(ins[33]), .en, .reset(rst), .clk);
	FF_en r32(.q(outs[32]), .d(ins[32]), .en, .reset(rst), .clk);
		FF_en r47(.q(outs[47]), .d(ins[47]), .en, .reset(rst), .clk);
	FF_en r46(.q(outs[46]), .d(ins[46]), .en, .reset(rst), .clk);
	FF_en r45(.q(outs[45]), .d(ins[45]), .en, .reset(rst), .clk);
	FF_en r44(.q(outs[44]), .d(ins[44]), .en, .reset(rst), .clk);
	FF_en r43(.q(outs[43]), .d(ins[43]), .en, .reset(rst), .clk);
	FF_en r42(.q(outs[42]), .d(ins[42]), .en, .reset(rst), .clk);
	FF_en r41(.q(outs[41]), .d(ins[41]), .en, .reset(rst), .clk);
	FF_en r40(.q(outs[40]), .d(ins[40]), .en, .reset(rst), .clk);
		FF_en r55(.q(outs[55]), .d(ins[55]), .en, .reset(rst), .clk);
	FF_en r54(.q(outs[54]), .d(ins[54]), .en, .reset(rst), .clk);
	FF_en r53(.q(outs[53]), .d(ins[53]), .en, .reset(rst), .clk);
	FF_en r52(.q(outs[52]), .d(ins[52]), .en, .reset(rst), .clk);
	FF_en r51(.q(outs[51]), .d(ins[51]), .en, .reset(rst), .clk);
	FF_en r50(.q(outs[50]), .d(ins[50]), .en, .reset(rst), .clk);
	FF_en r49(.q(outs[49]), .d(ins[49]), .en, .reset(rst), .clk);
	FF_en r48(.q(outs[48]), .d(ins[48]), .en, .reset(rst), .clk);
		FF_en r63(.q(outs[63]), .d(ins[63]), .en, .reset(rst), .clk);
	FF_en r62(.q(outs[62]), .d(ins[62]), .en, .reset(rst), .clk);
	FF_en r61(.q(outs[61]), .d(ins[61]), .en, .reset(rst), .clk);
	FF_en r60(.q(outs[60]), .d(ins[60]), .en, .reset(rst), .clk);
	FF_en r59(.q(outs[59]), .d(ins[59]), .en, .reset(rst), .clk);
	FF_en r58(.q(outs[58]), .d(ins[58]), .en, .reset(rst), .clk);
	FF_en r57(.q(outs[57]), .d(ins[57]), .en, .reset(rst), .clk);
	FF_en r56(.q(outs[56]), .d(ins[56]), .en, .reset(rst), .clk);
endmodule

